module \std::conv::bit_to_bool  (
        input b_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::bit_to_bool" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::bit_to_bool );
        end
    end
    `endif
    logic \b ;
    assign \b  = b_i;
    logic _e_1;
    assign _e_1 = \b ;
    assign output__ = _e_1;
endmodule

module \std::conv::unsafe::clock_to_bool  (
        input c_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::unsafe::clock_to_bool" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::unsafe::clock_to_bool );
        end
    end
    `endif
    logic \c ;
    assign \c  = c_i;
    logic _e_22;
    assign _e_22 = \c ;
    assign output__ = _e_22;
endmodule

module \std::conv::unsafe::bool_to_clock  (
        input c_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::unsafe::bool_to_clock" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::unsafe::bool_to_clock );
        end
    end
    `endif
    logic \c ;
    assign \c  = c_i;
    logic _e_25;
    assign _e_25 = \c ;
    assign output__ = _e_25;
endmodule

module \std::io::rising_edge  (
        input clk_i,
        input sync1_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::io::rising_edge" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::io::rising_edge );
        end
    end
    `endif
    logic \clk ;
    assign \clk  = clk_i;
    logic \sync1 ;
    assign \sync1  = sync1_i;
    (* src = "<compiler dir>/stdlib/io.spade:3,14" *)
    reg \sync2 ;
    (* src = "<compiler dir>/stdlib/io.spade:4,14" *)
    logic _e_33;
    (* src = "<compiler dir>/stdlib/io.spade:4,5" *)
    logic _e_31;
    always @(posedge \clk ) begin
        \sync2  <= \sync1 ;
    end
    assign _e_33 = !\sync2 ;
    assign _e_31 = \sync1  && _e_33;
    assign output__ = _e_31;
endmodule

module \std::io::falling_edge  (
        input clk_i,
        input sync1_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::io::falling_edge" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::io::falling_edge );
        end
    end
    `endif
    logic \clk ;
    assign \clk  = clk_i;
    logic \sync1 ;
    assign \sync1  = sync1_i;
    (* src = "<compiler dir>/stdlib/io.spade:9,14" *)
    reg \sync2 ;
    (* src = "<compiler dir>/stdlib/io.spade:10,14" *)
    logic _e_41;
    (* src = "<compiler dir>/stdlib/io.spade:10,5" *)
    logic _e_39;
    always @(posedge \clk ) begin
        \sync2  <= \sync1 ;
    end
    assign _e_41 = !\sync1 ;
    assign _e_39 = \sync2  && _e_41;
    assign output__ = _e_39;
endmodule

module \std::cdc::sync2_bool  (
        input clk_i,
        input in_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::cdc::sync2_bool" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::cdc::sync2_bool );
        end
    end
    `endif
    logic \clk ;
    assign \clk  = clk_i;
    logic \in ;
    assign \in  = in_i;
    (* src = "<compiler dir>/stdlib/cdc.spade:38,5" *)
    logic _e_335;
    (* src = "<compiler dir>/stdlib/cdc.spade:38,5" *)
    \std::cdc::unsafe::sync2[345]  sync2_0(.clk_i(\clk ), .in_i(\in ), .output__(_e_335));
    assign output__ = _e_335;
endmodule

module \tt07_delay_line_tmng::main::shift_reg  (
        input clk_i,
        input feedback_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "tt07_delay_line_tmng::main::shift_reg" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \tt07_delay_line_tmng::main::shift_reg );
        end
    end
    `endif
    logic \clk ;
    assign \clk  = clk_i;
    logic \feedback ;
    assign \feedback  = feedback_i;
    (* src = "src/main.spade:4,5" *)
    reg \s1_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s2_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s3_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s4_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s5_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s6_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s7_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s8_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s9_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s10_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s11_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s12_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s13_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s14_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s15_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s16_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s17_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s18_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s19_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s20_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s21_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s22_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s23_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s24_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s25_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s26_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s27_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s28_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s29_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s30_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s31_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s32_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s33_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s34_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s35_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s36_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s37_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s38_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s39_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s40_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s41_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s42_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s43_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s44_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s45_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s46_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s47_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s48_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s49_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s50_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s51_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s52_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s53_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s54_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s55_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s56_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s57_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s58_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s59_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s60_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s61_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s62_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s63_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s64_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s65_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s66_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s67_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s68_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s69_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s70_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s71_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s72_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s73_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s74_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s75_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s76_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s77_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s78_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s79_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s80_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s81_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s82_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s83_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s84_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s85_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s86_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s87_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s88_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s89_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s90_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s91_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s92_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s93_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s94_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s95_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s96_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s97_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s98_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s99_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s100_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s101_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s102_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s103_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s104_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s105_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s106_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s107_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s108_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s109_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s110_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s111_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s112_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s113_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s114_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s115_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s116_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s117_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s118_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s119_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s120_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s121_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s122_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s123_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s124_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s125_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s126_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s127_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s128_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s129_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s130_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s131_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s132_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s133_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s134_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s135_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s136_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s137_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s138_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s139_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s140_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s141_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s142_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s143_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s144_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s145_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s146_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s147_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s148_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s149_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s150_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s151_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s152_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s153_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s154_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s155_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s156_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s157_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s158_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s159_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s160_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s161_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s162_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s163_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s164_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s165_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s166_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s167_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s168_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s169_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s170_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s171_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s172_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s173_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s174_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s175_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s176_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s177_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s178_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s179_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s180_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s181_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s182_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s183_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s184_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s185_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s186_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s187_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s188_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s189_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s190_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s191_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s192_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s193_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s194_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s195_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s196_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s197_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s198_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s199_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s200_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s201_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s202_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s203_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s204_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s205_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s206_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s207_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s208_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s209_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s210_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s211_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s212_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s213_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s214_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s215_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s216_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s217_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s218_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s219_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s220_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s221_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s222_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s223_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s224_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s225_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s226_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s227_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s228_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s229_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s230_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s231_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s232_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s233_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s234_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s235_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s236_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s237_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s238_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s239_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s240_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s241_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s242_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s243_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s244_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s245_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s246_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s247_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s248_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s249_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s250_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s251_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s252_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s253_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s254_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s255_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s256_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s257_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s258_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s259_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s260_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s261_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s262_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s263_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s264_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s265_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s266_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s267_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s268_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s269_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s270_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s271_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s272_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s273_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s274_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s275_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s276_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s277_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s278_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s279_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s280_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s281_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s282_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s283_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s284_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s285_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s286_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s287_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s288_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s289_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s290_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s291_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s292_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s293_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s294_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s295_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s296_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s297_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s298_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s299_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s300_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s301_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s302_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s303_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s304_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s305_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s306_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s307_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s308_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s309_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s310_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s311_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s312_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s313_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s314_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s315_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s316_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s317_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s318_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s319_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s320_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s321_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s322_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s323_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s324_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s325_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s326_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s327_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s328_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s329_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s330_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s331_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s332_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s333_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s334_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s335_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s336_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s337_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s338_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s339_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s340_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s341_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s342_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s343_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s344_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s345_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s346_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s347_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s348_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s349_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s350_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s351_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s352_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s353_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s354_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s355_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s356_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s357_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s358_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s359_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s360_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s361_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s362_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s363_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s364_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s365_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s366_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s367_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s368_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s369_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s370_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s371_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s372_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s373_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s374_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s375_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s376_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s377_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s378_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s379_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s380_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s381_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s382_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s383_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s384_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s385_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s386_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s387_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s388_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s389_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s390_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s391_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s392_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s393_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s394_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s395_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s396_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s397_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s398_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s399_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s400_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s401_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s402_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s403_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s404_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s405_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s406_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s407_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s408_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s409_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s410_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s411_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s412_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s413_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s414_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s415_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s416_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s417_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s418_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s419_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s420_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s421_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s422_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s423_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s424_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s425_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s426_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s427_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s428_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s429_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s430_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s431_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s432_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s433_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s434_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s435_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s436_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s437_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s438_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s439_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s440_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s441_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s442_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s443_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s444_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s445_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s446_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s447_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s448_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s449_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s450_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s451_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s452_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s453_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s454_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s455_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s456_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s457_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s458_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s459_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s460_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s461_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s462_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s463_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s464_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s465_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s466_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s467_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s468_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s469_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s470_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s471_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s472_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s473_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s474_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s475_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s476_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s477_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s478_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s479_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s480_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s481_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s482_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s483_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s484_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s485_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s486_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s487_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s488_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s489_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s490_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s491_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s492_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s493_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s494_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s495_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s496_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s497_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s498_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s499_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s500_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s501_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s502_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s503_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s504_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s505_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s506_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s507_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s508_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s509_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s510_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s511_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s512_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s513_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s514_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s515_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s516_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s517_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s518_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s519_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s520_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s521_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s522_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s523_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s524_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s525_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s526_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s527_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s528_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s529_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s530_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s531_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s532_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s533_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s534_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s535_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s536_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s537_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s538_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s539_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s540_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s541_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s542_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s543_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s544_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s545_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s546_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s547_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s548_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s549_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s550_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s551_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s552_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s553_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s554_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s555_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s556_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s557_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s558_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s559_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s560_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s561_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s562_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s563_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s564_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s565_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s566_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s567_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s568_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s569_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s570_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s571_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s572_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s573_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s574_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s575_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s576_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s577_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s578_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s579_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s580_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s581_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s582_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s583_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s584_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s585_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s586_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s587_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s588_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s589_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s590_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s591_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s592_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s593_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s594_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s595_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s596_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s597_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s598_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s599_feedback ;
    (* src = "src/main.spade:4,5" *)
    reg \s600_feedback ;
    always @(posedge \clk ) begin
        \s1_feedback  <= \feedback ;
    end
    always @(posedge \clk ) begin
        \s2_feedback  <= \s1_feedback ;
    end
    always @(posedge \clk ) begin
        \s3_feedback  <= \s2_feedback ;
    end
    always @(posedge \clk ) begin
        \s4_feedback  <= \s3_feedback ;
    end
    always @(posedge \clk ) begin
        \s5_feedback  <= \s4_feedback ;
    end
    always @(posedge \clk ) begin
        \s6_feedback  <= \s5_feedback ;
    end
    always @(posedge \clk ) begin
        \s7_feedback  <= \s6_feedback ;
    end
    always @(posedge \clk ) begin
        \s8_feedback  <= \s7_feedback ;
    end
    always @(posedge \clk ) begin
        \s9_feedback  <= \s8_feedback ;
    end
    always @(posedge \clk ) begin
        \s10_feedback  <= \s9_feedback ;
    end
    always @(posedge \clk ) begin
        \s11_feedback  <= \s10_feedback ;
    end
    always @(posedge \clk ) begin
        \s12_feedback  <= \s11_feedback ;
    end
    always @(posedge \clk ) begin
        \s13_feedback  <= \s12_feedback ;
    end
    always @(posedge \clk ) begin
        \s14_feedback  <= \s13_feedback ;
    end
    always @(posedge \clk ) begin
        \s15_feedback  <= \s14_feedback ;
    end
    always @(posedge \clk ) begin
        \s16_feedback  <= \s15_feedback ;
    end
    always @(posedge \clk ) begin
        \s17_feedback  <= \s16_feedback ;
    end
    always @(posedge \clk ) begin
        \s18_feedback  <= \s17_feedback ;
    end
    always @(posedge \clk ) begin
        \s19_feedback  <= \s18_feedback ;
    end
    always @(posedge \clk ) begin
        \s20_feedback  <= \s19_feedback ;
    end
    always @(posedge \clk ) begin
        \s21_feedback  <= \s20_feedback ;
    end
    always @(posedge \clk ) begin
        \s22_feedback  <= \s21_feedback ;
    end
    always @(posedge \clk ) begin
        \s23_feedback  <= \s22_feedback ;
    end
    always @(posedge \clk ) begin
        \s24_feedback  <= \s23_feedback ;
    end
    always @(posedge \clk ) begin
        \s25_feedback  <= \s24_feedback ;
    end
    always @(posedge \clk ) begin
        \s26_feedback  <= \s25_feedback ;
    end
    always @(posedge \clk ) begin
        \s27_feedback  <= \s26_feedback ;
    end
    always @(posedge \clk ) begin
        \s28_feedback  <= \s27_feedback ;
    end
    always @(posedge \clk ) begin
        \s29_feedback  <= \s28_feedback ;
    end
    always @(posedge \clk ) begin
        \s30_feedback  <= \s29_feedback ;
    end
    always @(posedge \clk ) begin
        \s31_feedback  <= \s30_feedback ;
    end
    always @(posedge \clk ) begin
        \s32_feedback  <= \s31_feedback ;
    end
    always @(posedge \clk ) begin
        \s33_feedback  <= \s32_feedback ;
    end
    always @(posedge \clk ) begin
        \s34_feedback  <= \s33_feedback ;
    end
    always @(posedge \clk ) begin
        \s35_feedback  <= \s34_feedback ;
    end
    always @(posedge \clk ) begin
        \s36_feedback  <= \s35_feedback ;
    end
    always @(posedge \clk ) begin
        \s37_feedback  <= \s36_feedback ;
    end
    always @(posedge \clk ) begin
        \s38_feedback  <= \s37_feedback ;
    end
    always @(posedge \clk ) begin
        \s39_feedback  <= \s38_feedback ;
    end
    always @(posedge \clk ) begin
        \s40_feedback  <= \s39_feedback ;
    end
    always @(posedge \clk ) begin
        \s41_feedback  <= \s40_feedback ;
    end
    always @(posedge \clk ) begin
        \s42_feedback  <= \s41_feedback ;
    end
    always @(posedge \clk ) begin
        \s43_feedback  <= \s42_feedback ;
    end
    always @(posedge \clk ) begin
        \s44_feedback  <= \s43_feedback ;
    end
    always @(posedge \clk ) begin
        \s45_feedback  <= \s44_feedback ;
    end
    always @(posedge \clk ) begin
        \s46_feedback  <= \s45_feedback ;
    end
    always @(posedge \clk ) begin
        \s47_feedback  <= \s46_feedback ;
    end
    always @(posedge \clk ) begin
        \s48_feedback  <= \s47_feedback ;
    end
    always @(posedge \clk ) begin
        \s49_feedback  <= \s48_feedback ;
    end
    always @(posedge \clk ) begin
        \s50_feedback  <= \s49_feedback ;
    end
    always @(posedge \clk ) begin
        \s51_feedback  <= \s50_feedback ;
    end
    always @(posedge \clk ) begin
        \s52_feedback  <= \s51_feedback ;
    end
    always @(posedge \clk ) begin
        \s53_feedback  <= \s52_feedback ;
    end
    always @(posedge \clk ) begin
        \s54_feedback  <= \s53_feedback ;
    end
    always @(posedge \clk ) begin
        \s55_feedback  <= \s54_feedback ;
    end
    always @(posedge \clk ) begin
        \s56_feedback  <= \s55_feedback ;
    end
    always @(posedge \clk ) begin
        \s57_feedback  <= \s56_feedback ;
    end
    always @(posedge \clk ) begin
        \s58_feedback  <= \s57_feedback ;
    end
    always @(posedge \clk ) begin
        \s59_feedback  <= \s58_feedback ;
    end
    always @(posedge \clk ) begin
        \s60_feedback  <= \s59_feedback ;
    end
    always @(posedge \clk ) begin
        \s61_feedback  <= \s60_feedback ;
    end
    always @(posedge \clk ) begin
        \s62_feedback  <= \s61_feedback ;
    end
    always @(posedge \clk ) begin
        \s63_feedback  <= \s62_feedback ;
    end
    always @(posedge \clk ) begin
        \s64_feedback  <= \s63_feedback ;
    end
    always @(posedge \clk ) begin
        \s65_feedback  <= \s64_feedback ;
    end
    always @(posedge \clk ) begin
        \s66_feedback  <= \s65_feedback ;
    end
    always @(posedge \clk ) begin
        \s67_feedback  <= \s66_feedback ;
    end
    always @(posedge \clk ) begin
        \s68_feedback  <= \s67_feedback ;
    end
    always @(posedge \clk ) begin
        \s69_feedback  <= \s68_feedback ;
    end
    always @(posedge \clk ) begin
        \s70_feedback  <= \s69_feedback ;
    end
    always @(posedge \clk ) begin
        \s71_feedback  <= \s70_feedback ;
    end
    always @(posedge \clk ) begin
        \s72_feedback  <= \s71_feedback ;
    end
    always @(posedge \clk ) begin
        \s73_feedback  <= \s72_feedback ;
    end
    always @(posedge \clk ) begin
        \s74_feedback  <= \s73_feedback ;
    end
    always @(posedge \clk ) begin
        \s75_feedback  <= \s74_feedback ;
    end
    always @(posedge \clk ) begin
        \s76_feedback  <= \s75_feedback ;
    end
    always @(posedge \clk ) begin
        \s77_feedback  <= \s76_feedback ;
    end
    always @(posedge \clk ) begin
        \s78_feedback  <= \s77_feedback ;
    end
    always @(posedge \clk ) begin
        \s79_feedback  <= \s78_feedback ;
    end
    always @(posedge \clk ) begin
        \s80_feedback  <= \s79_feedback ;
    end
    always @(posedge \clk ) begin
        \s81_feedback  <= \s80_feedback ;
    end
    always @(posedge \clk ) begin
        \s82_feedback  <= \s81_feedback ;
    end
    always @(posedge \clk ) begin
        \s83_feedback  <= \s82_feedback ;
    end
    always @(posedge \clk ) begin
        \s84_feedback  <= \s83_feedback ;
    end
    always @(posedge \clk ) begin
        \s85_feedback  <= \s84_feedback ;
    end
    always @(posedge \clk ) begin
        \s86_feedback  <= \s85_feedback ;
    end
    always @(posedge \clk ) begin
        \s87_feedback  <= \s86_feedback ;
    end
    always @(posedge \clk ) begin
        \s88_feedback  <= \s87_feedback ;
    end
    always @(posedge \clk ) begin
        \s89_feedback  <= \s88_feedback ;
    end
    always @(posedge \clk ) begin
        \s90_feedback  <= \s89_feedback ;
    end
    always @(posedge \clk ) begin
        \s91_feedback  <= \s90_feedback ;
    end
    always @(posedge \clk ) begin
        \s92_feedback  <= \s91_feedback ;
    end
    always @(posedge \clk ) begin
        \s93_feedback  <= \s92_feedback ;
    end
    always @(posedge \clk ) begin
        \s94_feedback  <= \s93_feedback ;
    end
    always @(posedge \clk ) begin
        \s95_feedback  <= \s94_feedback ;
    end
    always @(posedge \clk ) begin
        \s96_feedback  <= \s95_feedback ;
    end
    always @(posedge \clk ) begin
        \s97_feedback  <= \s96_feedback ;
    end
    always @(posedge \clk ) begin
        \s98_feedback  <= \s97_feedback ;
    end
    always @(posedge \clk ) begin
        \s99_feedback  <= \s98_feedback ;
    end
    always @(posedge \clk ) begin
        \s100_feedback  <= \s99_feedback ;
    end
    always @(posedge \clk ) begin
        \s101_feedback  <= \s100_feedback ;
    end
    always @(posedge \clk ) begin
        \s102_feedback  <= \s101_feedback ;
    end
    always @(posedge \clk ) begin
        \s103_feedback  <= \s102_feedback ;
    end
    always @(posedge \clk ) begin
        \s104_feedback  <= \s103_feedback ;
    end
    always @(posedge \clk ) begin
        \s105_feedback  <= \s104_feedback ;
    end
    always @(posedge \clk ) begin
        \s106_feedback  <= \s105_feedback ;
    end
    always @(posedge \clk ) begin
        \s107_feedback  <= \s106_feedback ;
    end
    always @(posedge \clk ) begin
        \s108_feedback  <= \s107_feedback ;
    end
    always @(posedge \clk ) begin
        \s109_feedback  <= \s108_feedback ;
    end
    always @(posedge \clk ) begin
        \s110_feedback  <= \s109_feedback ;
    end
    always @(posedge \clk ) begin
        \s111_feedback  <= \s110_feedback ;
    end
    always @(posedge \clk ) begin
        \s112_feedback  <= \s111_feedback ;
    end
    always @(posedge \clk ) begin
        \s113_feedback  <= \s112_feedback ;
    end
    always @(posedge \clk ) begin
        \s114_feedback  <= \s113_feedback ;
    end
    always @(posedge \clk ) begin
        \s115_feedback  <= \s114_feedback ;
    end
    always @(posedge \clk ) begin
        \s116_feedback  <= \s115_feedback ;
    end
    always @(posedge \clk ) begin
        \s117_feedback  <= \s116_feedback ;
    end
    always @(posedge \clk ) begin
        \s118_feedback  <= \s117_feedback ;
    end
    always @(posedge \clk ) begin
        \s119_feedback  <= \s118_feedback ;
    end
    always @(posedge \clk ) begin
        \s120_feedback  <= \s119_feedback ;
    end
    always @(posedge \clk ) begin
        \s121_feedback  <= \s120_feedback ;
    end
    always @(posedge \clk ) begin
        \s122_feedback  <= \s121_feedback ;
    end
    always @(posedge \clk ) begin
        \s123_feedback  <= \s122_feedback ;
    end
    always @(posedge \clk ) begin
        \s124_feedback  <= \s123_feedback ;
    end
    always @(posedge \clk ) begin
        \s125_feedback  <= \s124_feedback ;
    end
    always @(posedge \clk ) begin
        \s126_feedback  <= \s125_feedback ;
    end
    always @(posedge \clk ) begin
        \s127_feedback  <= \s126_feedback ;
    end
    always @(posedge \clk ) begin
        \s128_feedback  <= \s127_feedback ;
    end
    always @(posedge \clk ) begin
        \s129_feedback  <= \s128_feedback ;
    end
    always @(posedge \clk ) begin
        \s130_feedback  <= \s129_feedback ;
    end
    always @(posedge \clk ) begin
        \s131_feedback  <= \s130_feedback ;
    end
    always @(posedge \clk ) begin
        \s132_feedback  <= \s131_feedback ;
    end
    always @(posedge \clk ) begin
        \s133_feedback  <= \s132_feedback ;
    end
    always @(posedge \clk ) begin
        \s134_feedback  <= \s133_feedback ;
    end
    always @(posedge \clk ) begin
        \s135_feedback  <= \s134_feedback ;
    end
    always @(posedge \clk ) begin
        \s136_feedback  <= \s135_feedback ;
    end
    always @(posedge \clk ) begin
        \s137_feedback  <= \s136_feedback ;
    end
    always @(posedge \clk ) begin
        \s138_feedback  <= \s137_feedback ;
    end
    always @(posedge \clk ) begin
        \s139_feedback  <= \s138_feedback ;
    end
    always @(posedge \clk ) begin
        \s140_feedback  <= \s139_feedback ;
    end
    always @(posedge \clk ) begin
        \s141_feedback  <= \s140_feedback ;
    end
    always @(posedge \clk ) begin
        \s142_feedback  <= \s141_feedback ;
    end
    always @(posedge \clk ) begin
        \s143_feedback  <= \s142_feedback ;
    end
    always @(posedge \clk ) begin
        \s144_feedback  <= \s143_feedback ;
    end
    always @(posedge \clk ) begin
        \s145_feedback  <= \s144_feedback ;
    end
    always @(posedge \clk ) begin
        \s146_feedback  <= \s145_feedback ;
    end
    always @(posedge \clk ) begin
        \s147_feedback  <= \s146_feedback ;
    end
    always @(posedge \clk ) begin
        \s148_feedback  <= \s147_feedback ;
    end
    always @(posedge \clk ) begin
        \s149_feedback  <= \s148_feedback ;
    end
    always @(posedge \clk ) begin
        \s150_feedback  <= \s149_feedback ;
    end
    always @(posedge \clk ) begin
        \s151_feedback  <= \s150_feedback ;
    end
    always @(posedge \clk ) begin
        \s152_feedback  <= \s151_feedback ;
    end
    always @(posedge \clk ) begin
        \s153_feedback  <= \s152_feedback ;
    end
    always @(posedge \clk ) begin
        \s154_feedback  <= \s153_feedback ;
    end
    always @(posedge \clk ) begin
        \s155_feedback  <= \s154_feedback ;
    end
    always @(posedge \clk ) begin
        \s156_feedback  <= \s155_feedback ;
    end
    always @(posedge \clk ) begin
        \s157_feedback  <= \s156_feedback ;
    end
    always @(posedge \clk ) begin
        \s158_feedback  <= \s157_feedback ;
    end
    always @(posedge \clk ) begin
        \s159_feedback  <= \s158_feedback ;
    end
    always @(posedge \clk ) begin
        \s160_feedback  <= \s159_feedback ;
    end
    always @(posedge \clk ) begin
        \s161_feedback  <= \s160_feedback ;
    end
    always @(posedge \clk ) begin
        \s162_feedback  <= \s161_feedback ;
    end
    always @(posedge \clk ) begin
        \s163_feedback  <= \s162_feedback ;
    end
    always @(posedge \clk ) begin
        \s164_feedback  <= \s163_feedback ;
    end
    always @(posedge \clk ) begin
        \s165_feedback  <= \s164_feedback ;
    end
    always @(posedge \clk ) begin
        \s166_feedback  <= \s165_feedback ;
    end
    always @(posedge \clk ) begin
        \s167_feedback  <= \s166_feedback ;
    end
    always @(posedge \clk ) begin
        \s168_feedback  <= \s167_feedback ;
    end
    always @(posedge \clk ) begin
        \s169_feedback  <= \s168_feedback ;
    end
    always @(posedge \clk ) begin
        \s170_feedback  <= \s169_feedback ;
    end
    always @(posedge \clk ) begin
        \s171_feedback  <= \s170_feedback ;
    end
    always @(posedge \clk ) begin
        \s172_feedback  <= \s171_feedback ;
    end
    always @(posedge \clk ) begin
        \s173_feedback  <= \s172_feedback ;
    end
    always @(posedge \clk ) begin
        \s174_feedback  <= \s173_feedback ;
    end
    always @(posedge \clk ) begin
        \s175_feedback  <= \s174_feedback ;
    end
    always @(posedge \clk ) begin
        \s176_feedback  <= \s175_feedback ;
    end
    always @(posedge \clk ) begin
        \s177_feedback  <= \s176_feedback ;
    end
    always @(posedge \clk ) begin
        \s178_feedback  <= \s177_feedback ;
    end
    always @(posedge \clk ) begin
        \s179_feedback  <= \s178_feedback ;
    end
    always @(posedge \clk ) begin
        \s180_feedback  <= \s179_feedback ;
    end
    always @(posedge \clk ) begin
        \s181_feedback  <= \s180_feedback ;
    end
    always @(posedge \clk ) begin
        \s182_feedback  <= \s181_feedback ;
    end
    always @(posedge \clk ) begin
        \s183_feedback  <= \s182_feedback ;
    end
    always @(posedge \clk ) begin
        \s184_feedback  <= \s183_feedback ;
    end
    always @(posedge \clk ) begin
        \s185_feedback  <= \s184_feedback ;
    end
    always @(posedge \clk ) begin
        \s186_feedback  <= \s185_feedback ;
    end
    always @(posedge \clk ) begin
        \s187_feedback  <= \s186_feedback ;
    end
    always @(posedge \clk ) begin
        \s188_feedback  <= \s187_feedback ;
    end
    always @(posedge \clk ) begin
        \s189_feedback  <= \s188_feedback ;
    end
    always @(posedge \clk ) begin
        \s190_feedback  <= \s189_feedback ;
    end
    always @(posedge \clk ) begin
        \s191_feedback  <= \s190_feedback ;
    end
    always @(posedge \clk ) begin
        \s192_feedback  <= \s191_feedback ;
    end
    always @(posedge \clk ) begin
        \s193_feedback  <= \s192_feedback ;
    end
    always @(posedge \clk ) begin
        \s194_feedback  <= \s193_feedback ;
    end
    always @(posedge \clk ) begin
        \s195_feedback  <= \s194_feedback ;
    end
    always @(posedge \clk ) begin
        \s196_feedback  <= \s195_feedback ;
    end
    always @(posedge \clk ) begin
        \s197_feedback  <= \s196_feedback ;
    end
    always @(posedge \clk ) begin
        \s198_feedback  <= \s197_feedback ;
    end
    always @(posedge \clk ) begin
        \s199_feedback  <= \s198_feedback ;
    end
    always @(posedge \clk ) begin
        \s200_feedback  <= \s199_feedback ;
    end
    always @(posedge \clk ) begin
        \s201_feedback  <= \s200_feedback ;
    end
    always @(posedge \clk ) begin
        \s202_feedback  <= \s201_feedback ;
    end
    always @(posedge \clk ) begin
        \s203_feedback  <= \s202_feedback ;
    end
    always @(posedge \clk ) begin
        \s204_feedback  <= \s203_feedback ;
    end
    always @(posedge \clk ) begin
        \s205_feedback  <= \s204_feedback ;
    end
    always @(posedge \clk ) begin
        \s206_feedback  <= \s205_feedback ;
    end
    always @(posedge \clk ) begin
        \s207_feedback  <= \s206_feedback ;
    end
    always @(posedge \clk ) begin
        \s208_feedback  <= \s207_feedback ;
    end
    always @(posedge \clk ) begin
        \s209_feedback  <= \s208_feedback ;
    end
    always @(posedge \clk ) begin
        \s210_feedback  <= \s209_feedback ;
    end
    always @(posedge \clk ) begin
        \s211_feedback  <= \s210_feedback ;
    end
    always @(posedge \clk ) begin
        \s212_feedback  <= \s211_feedback ;
    end
    always @(posedge \clk ) begin
        \s213_feedback  <= \s212_feedback ;
    end
    always @(posedge \clk ) begin
        \s214_feedback  <= \s213_feedback ;
    end
    always @(posedge \clk ) begin
        \s215_feedback  <= \s214_feedback ;
    end
    always @(posedge \clk ) begin
        \s216_feedback  <= \s215_feedback ;
    end
    always @(posedge \clk ) begin
        \s217_feedback  <= \s216_feedback ;
    end
    always @(posedge \clk ) begin
        \s218_feedback  <= \s217_feedback ;
    end
    always @(posedge \clk ) begin
        \s219_feedback  <= \s218_feedback ;
    end
    always @(posedge \clk ) begin
        \s220_feedback  <= \s219_feedback ;
    end
    always @(posedge \clk ) begin
        \s221_feedback  <= \s220_feedback ;
    end
    always @(posedge \clk ) begin
        \s222_feedback  <= \s221_feedback ;
    end
    always @(posedge \clk ) begin
        \s223_feedback  <= \s222_feedback ;
    end
    always @(posedge \clk ) begin
        \s224_feedback  <= \s223_feedback ;
    end
    always @(posedge \clk ) begin
        \s225_feedback  <= \s224_feedback ;
    end
    always @(posedge \clk ) begin
        \s226_feedback  <= \s225_feedback ;
    end
    always @(posedge \clk ) begin
        \s227_feedback  <= \s226_feedback ;
    end
    always @(posedge \clk ) begin
        \s228_feedback  <= \s227_feedback ;
    end
    always @(posedge \clk ) begin
        \s229_feedback  <= \s228_feedback ;
    end
    always @(posedge \clk ) begin
        \s230_feedback  <= \s229_feedback ;
    end
    always @(posedge \clk ) begin
        \s231_feedback  <= \s230_feedback ;
    end
    always @(posedge \clk ) begin
        \s232_feedback  <= \s231_feedback ;
    end
    always @(posedge \clk ) begin
        \s233_feedback  <= \s232_feedback ;
    end
    always @(posedge \clk ) begin
        \s234_feedback  <= \s233_feedback ;
    end
    always @(posedge \clk ) begin
        \s235_feedback  <= \s234_feedback ;
    end
    always @(posedge \clk ) begin
        \s236_feedback  <= \s235_feedback ;
    end
    always @(posedge \clk ) begin
        \s237_feedback  <= \s236_feedback ;
    end
    always @(posedge \clk ) begin
        \s238_feedback  <= \s237_feedback ;
    end
    always @(posedge \clk ) begin
        \s239_feedback  <= \s238_feedback ;
    end
    always @(posedge \clk ) begin
        \s240_feedback  <= \s239_feedback ;
    end
    always @(posedge \clk ) begin
        \s241_feedback  <= \s240_feedback ;
    end
    always @(posedge \clk ) begin
        \s242_feedback  <= \s241_feedback ;
    end
    always @(posedge \clk ) begin
        \s243_feedback  <= \s242_feedback ;
    end
    always @(posedge \clk ) begin
        \s244_feedback  <= \s243_feedback ;
    end
    always @(posedge \clk ) begin
        \s245_feedback  <= \s244_feedback ;
    end
    always @(posedge \clk ) begin
        \s246_feedback  <= \s245_feedback ;
    end
    always @(posedge \clk ) begin
        \s247_feedback  <= \s246_feedback ;
    end
    always @(posedge \clk ) begin
        \s248_feedback  <= \s247_feedback ;
    end
    always @(posedge \clk ) begin
        \s249_feedback  <= \s248_feedback ;
    end
    always @(posedge \clk ) begin
        \s250_feedback  <= \s249_feedback ;
    end
    always @(posedge \clk ) begin
        \s251_feedback  <= \s250_feedback ;
    end
    always @(posedge \clk ) begin
        \s252_feedback  <= \s251_feedback ;
    end
    always @(posedge \clk ) begin
        \s253_feedback  <= \s252_feedback ;
    end
    always @(posedge \clk ) begin
        \s254_feedback  <= \s253_feedback ;
    end
    always @(posedge \clk ) begin
        \s255_feedback  <= \s254_feedback ;
    end
    always @(posedge \clk ) begin
        \s256_feedback  <= \s255_feedback ;
    end
    always @(posedge \clk ) begin
        \s257_feedback  <= \s256_feedback ;
    end
    always @(posedge \clk ) begin
        \s258_feedback  <= \s257_feedback ;
    end
    always @(posedge \clk ) begin
        \s259_feedback  <= \s258_feedback ;
    end
    always @(posedge \clk ) begin
        \s260_feedback  <= \s259_feedback ;
    end
    always @(posedge \clk ) begin
        \s261_feedback  <= \s260_feedback ;
    end
    always @(posedge \clk ) begin
        \s262_feedback  <= \s261_feedback ;
    end
    always @(posedge \clk ) begin
        \s263_feedback  <= \s262_feedback ;
    end
    always @(posedge \clk ) begin
        \s264_feedback  <= \s263_feedback ;
    end
    always @(posedge \clk ) begin
        \s265_feedback  <= \s264_feedback ;
    end
    always @(posedge \clk ) begin
        \s266_feedback  <= \s265_feedback ;
    end
    always @(posedge \clk ) begin
        \s267_feedback  <= \s266_feedback ;
    end
    always @(posedge \clk ) begin
        \s268_feedback  <= \s267_feedback ;
    end
    always @(posedge \clk ) begin
        \s269_feedback  <= \s268_feedback ;
    end
    always @(posedge \clk ) begin
        \s270_feedback  <= \s269_feedback ;
    end
    always @(posedge \clk ) begin
        \s271_feedback  <= \s270_feedback ;
    end
    always @(posedge \clk ) begin
        \s272_feedback  <= \s271_feedback ;
    end
    always @(posedge \clk ) begin
        \s273_feedback  <= \s272_feedback ;
    end
    always @(posedge \clk ) begin
        \s274_feedback  <= \s273_feedback ;
    end
    always @(posedge \clk ) begin
        \s275_feedback  <= \s274_feedback ;
    end
    always @(posedge \clk ) begin
        \s276_feedback  <= \s275_feedback ;
    end
    always @(posedge \clk ) begin
        \s277_feedback  <= \s276_feedback ;
    end
    always @(posedge \clk ) begin
        \s278_feedback  <= \s277_feedback ;
    end
    always @(posedge \clk ) begin
        \s279_feedback  <= \s278_feedback ;
    end
    always @(posedge \clk ) begin
        \s280_feedback  <= \s279_feedback ;
    end
    always @(posedge \clk ) begin
        \s281_feedback  <= \s280_feedback ;
    end
    always @(posedge \clk ) begin
        \s282_feedback  <= \s281_feedback ;
    end
    always @(posedge \clk ) begin
        \s283_feedback  <= \s282_feedback ;
    end
    always @(posedge \clk ) begin
        \s284_feedback  <= \s283_feedback ;
    end
    always @(posedge \clk ) begin
        \s285_feedback  <= \s284_feedback ;
    end
    always @(posedge \clk ) begin
        \s286_feedback  <= \s285_feedback ;
    end
    always @(posedge \clk ) begin
        \s287_feedback  <= \s286_feedback ;
    end
    always @(posedge \clk ) begin
        \s288_feedback  <= \s287_feedback ;
    end
    always @(posedge \clk ) begin
        \s289_feedback  <= \s288_feedback ;
    end
    always @(posedge \clk ) begin
        \s290_feedback  <= \s289_feedback ;
    end
    always @(posedge \clk ) begin
        \s291_feedback  <= \s290_feedback ;
    end
    always @(posedge \clk ) begin
        \s292_feedback  <= \s291_feedback ;
    end
    always @(posedge \clk ) begin
        \s293_feedback  <= \s292_feedback ;
    end
    always @(posedge \clk ) begin
        \s294_feedback  <= \s293_feedback ;
    end
    always @(posedge \clk ) begin
        \s295_feedback  <= \s294_feedback ;
    end
    always @(posedge \clk ) begin
        \s296_feedback  <= \s295_feedback ;
    end
    always @(posedge \clk ) begin
        \s297_feedback  <= \s296_feedback ;
    end
    always @(posedge \clk ) begin
        \s298_feedback  <= \s297_feedback ;
    end
    always @(posedge \clk ) begin
        \s299_feedback  <= \s298_feedback ;
    end
    always @(posedge \clk ) begin
        \s300_feedback  <= \s299_feedback ;
    end
    always @(posedge \clk ) begin
        \s301_feedback  <= \s300_feedback ;
    end
    always @(posedge \clk ) begin
        \s302_feedback  <= \s301_feedback ;
    end
    always @(posedge \clk ) begin
        \s303_feedback  <= \s302_feedback ;
    end
    always @(posedge \clk ) begin
        \s304_feedback  <= \s303_feedback ;
    end
    always @(posedge \clk ) begin
        \s305_feedback  <= \s304_feedback ;
    end
    always @(posedge \clk ) begin
        \s306_feedback  <= \s305_feedback ;
    end
    always @(posedge \clk ) begin
        \s307_feedback  <= \s306_feedback ;
    end
    always @(posedge \clk ) begin
        \s308_feedback  <= \s307_feedback ;
    end
    always @(posedge \clk ) begin
        \s309_feedback  <= \s308_feedback ;
    end
    always @(posedge \clk ) begin
        \s310_feedback  <= \s309_feedback ;
    end
    always @(posedge \clk ) begin
        \s311_feedback  <= \s310_feedback ;
    end
    always @(posedge \clk ) begin
        \s312_feedback  <= \s311_feedback ;
    end
    always @(posedge \clk ) begin
        \s313_feedback  <= \s312_feedback ;
    end
    always @(posedge \clk ) begin
        \s314_feedback  <= \s313_feedback ;
    end
    always @(posedge \clk ) begin
        \s315_feedback  <= \s314_feedback ;
    end
    always @(posedge \clk ) begin
        \s316_feedback  <= \s315_feedback ;
    end
    always @(posedge \clk ) begin
        \s317_feedback  <= \s316_feedback ;
    end
    always @(posedge \clk ) begin
        \s318_feedback  <= \s317_feedback ;
    end
    always @(posedge \clk ) begin
        \s319_feedback  <= \s318_feedback ;
    end
    always @(posedge \clk ) begin
        \s320_feedback  <= \s319_feedback ;
    end
    always @(posedge \clk ) begin
        \s321_feedback  <= \s320_feedback ;
    end
    always @(posedge \clk ) begin
        \s322_feedback  <= \s321_feedback ;
    end
    always @(posedge \clk ) begin
        \s323_feedback  <= \s322_feedback ;
    end
    always @(posedge \clk ) begin
        \s324_feedback  <= \s323_feedback ;
    end
    always @(posedge \clk ) begin
        \s325_feedback  <= \s324_feedback ;
    end
    always @(posedge \clk ) begin
        \s326_feedback  <= \s325_feedback ;
    end
    always @(posedge \clk ) begin
        \s327_feedback  <= \s326_feedback ;
    end
    always @(posedge \clk ) begin
        \s328_feedback  <= \s327_feedback ;
    end
    always @(posedge \clk ) begin
        \s329_feedback  <= \s328_feedback ;
    end
    always @(posedge \clk ) begin
        \s330_feedback  <= \s329_feedback ;
    end
    always @(posedge \clk ) begin
        \s331_feedback  <= \s330_feedback ;
    end
    always @(posedge \clk ) begin
        \s332_feedback  <= \s331_feedback ;
    end
    always @(posedge \clk ) begin
        \s333_feedback  <= \s332_feedback ;
    end
    always @(posedge \clk ) begin
        \s334_feedback  <= \s333_feedback ;
    end
    always @(posedge \clk ) begin
        \s335_feedback  <= \s334_feedback ;
    end
    always @(posedge \clk ) begin
        \s336_feedback  <= \s335_feedback ;
    end
    always @(posedge \clk ) begin
        \s337_feedback  <= \s336_feedback ;
    end
    always @(posedge \clk ) begin
        \s338_feedback  <= \s337_feedback ;
    end
    always @(posedge \clk ) begin
        \s339_feedback  <= \s338_feedback ;
    end
    always @(posedge \clk ) begin
        \s340_feedback  <= \s339_feedback ;
    end
    always @(posedge \clk ) begin
        \s341_feedback  <= \s340_feedback ;
    end
    always @(posedge \clk ) begin
        \s342_feedback  <= \s341_feedback ;
    end
    always @(posedge \clk ) begin
        \s343_feedback  <= \s342_feedback ;
    end
    always @(posedge \clk ) begin
        \s344_feedback  <= \s343_feedback ;
    end
    always @(posedge \clk ) begin
        \s345_feedback  <= \s344_feedback ;
    end
    always @(posedge \clk ) begin
        \s346_feedback  <= \s345_feedback ;
    end
    always @(posedge \clk ) begin
        \s347_feedback  <= \s346_feedback ;
    end
    always @(posedge \clk ) begin
        \s348_feedback  <= \s347_feedback ;
    end
    always @(posedge \clk ) begin
        \s349_feedback  <= \s348_feedback ;
    end
    always @(posedge \clk ) begin
        \s350_feedback  <= \s349_feedback ;
    end
    always @(posedge \clk ) begin
        \s351_feedback  <= \s350_feedback ;
    end
    always @(posedge \clk ) begin
        \s352_feedback  <= \s351_feedback ;
    end
    always @(posedge \clk ) begin
        \s353_feedback  <= \s352_feedback ;
    end
    always @(posedge \clk ) begin
        \s354_feedback  <= \s353_feedback ;
    end
    always @(posedge \clk ) begin
        \s355_feedback  <= \s354_feedback ;
    end
    always @(posedge \clk ) begin
        \s356_feedback  <= \s355_feedback ;
    end
    always @(posedge \clk ) begin
        \s357_feedback  <= \s356_feedback ;
    end
    always @(posedge \clk ) begin
        \s358_feedback  <= \s357_feedback ;
    end
    always @(posedge \clk ) begin
        \s359_feedback  <= \s358_feedback ;
    end
    always @(posedge \clk ) begin
        \s360_feedback  <= \s359_feedback ;
    end
    always @(posedge \clk ) begin
        \s361_feedback  <= \s360_feedback ;
    end
    always @(posedge \clk ) begin
        \s362_feedback  <= \s361_feedback ;
    end
    always @(posedge \clk ) begin
        \s363_feedback  <= \s362_feedback ;
    end
    always @(posedge \clk ) begin
        \s364_feedback  <= \s363_feedback ;
    end
    always @(posedge \clk ) begin
        \s365_feedback  <= \s364_feedback ;
    end
    always @(posedge \clk ) begin
        \s366_feedback  <= \s365_feedback ;
    end
    always @(posedge \clk ) begin
        \s367_feedback  <= \s366_feedback ;
    end
    always @(posedge \clk ) begin
        \s368_feedback  <= \s367_feedback ;
    end
    always @(posedge \clk ) begin
        \s369_feedback  <= \s368_feedback ;
    end
    always @(posedge \clk ) begin
        \s370_feedback  <= \s369_feedback ;
    end
    always @(posedge \clk ) begin
        \s371_feedback  <= \s370_feedback ;
    end
    always @(posedge \clk ) begin
        \s372_feedback  <= \s371_feedback ;
    end
    always @(posedge \clk ) begin
        \s373_feedback  <= \s372_feedback ;
    end
    always @(posedge \clk ) begin
        \s374_feedback  <= \s373_feedback ;
    end
    always @(posedge \clk ) begin
        \s375_feedback  <= \s374_feedback ;
    end
    always @(posedge \clk ) begin
        \s376_feedback  <= \s375_feedback ;
    end
    always @(posedge \clk ) begin
        \s377_feedback  <= \s376_feedback ;
    end
    always @(posedge \clk ) begin
        \s378_feedback  <= \s377_feedback ;
    end
    always @(posedge \clk ) begin
        \s379_feedback  <= \s378_feedback ;
    end
    always @(posedge \clk ) begin
        \s380_feedback  <= \s379_feedback ;
    end
    always @(posedge \clk ) begin
        \s381_feedback  <= \s380_feedback ;
    end
    always @(posedge \clk ) begin
        \s382_feedback  <= \s381_feedback ;
    end
    always @(posedge \clk ) begin
        \s383_feedback  <= \s382_feedback ;
    end
    always @(posedge \clk ) begin
        \s384_feedback  <= \s383_feedback ;
    end
    always @(posedge \clk ) begin
        \s385_feedback  <= \s384_feedback ;
    end
    always @(posedge \clk ) begin
        \s386_feedback  <= \s385_feedback ;
    end
    always @(posedge \clk ) begin
        \s387_feedback  <= \s386_feedback ;
    end
    always @(posedge \clk ) begin
        \s388_feedback  <= \s387_feedback ;
    end
    always @(posedge \clk ) begin
        \s389_feedback  <= \s388_feedback ;
    end
    always @(posedge \clk ) begin
        \s390_feedback  <= \s389_feedback ;
    end
    always @(posedge \clk ) begin
        \s391_feedback  <= \s390_feedback ;
    end
    always @(posedge \clk ) begin
        \s392_feedback  <= \s391_feedback ;
    end
    always @(posedge \clk ) begin
        \s393_feedback  <= \s392_feedback ;
    end
    always @(posedge \clk ) begin
        \s394_feedback  <= \s393_feedback ;
    end
    always @(posedge \clk ) begin
        \s395_feedback  <= \s394_feedback ;
    end
    always @(posedge \clk ) begin
        \s396_feedback  <= \s395_feedback ;
    end
    always @(posedge \clk ) begin
        \s397_feedback  <= \s396_feedback ;
    end
    always @(posedge \clk ) begin
        \s398_feedback  <= \s397_feedback ;
    end
    always @(posedge \clk ) begin
        \s399_feedback  <= \s398_feedback ;
    end
    always @(posedge \clk ) begin
        \s400_feedback  <= \s399_feedback ;
    end
    always @(posedge \clk ) begin
        \s401_feedback  <= \s400_feedback ;
    end
    always @(posedge \clk ) begin
        \s402_feedback  <= \s401_feedback ;
    end
    always @(posedge \clk ) begin
        \s403_feedback  <= \s402_feedback ;
    end
    always @(posedge \clk ) begin
        \s404_feedback  <= \s403_feedback ;
    end
    always @(posedge \clk ) begin
        \s405_feedback  <= \s404_feedback ;
    end
    always @(posedge \clk ) begin
        \s406_feedback  <= \s405_feedback ;
    end
    always @(posedge \clk ) begin
        \s407_feedback  <= \s406_feedback ;
    end
    always @(posedge \clk ) begin
        \s408_feedback  <= \s407_feedback ;
    end
    always @(posedge \clk ) begin
        \s409_feedback  <= \s408_feedback ;
    end
    always @(posedge \clk ) begin
        \s410_feedback  <= \s409_feedback ;
    end
    always @(posedge \clk ) begin
        \s411_feedback  <= \s410_feedback ;
    end
    always @(posedge \clk ) begin
        \s412_feedback  <= \s411_feedback ;
    end
    always @(posedge \clk ) begin
        \s413_feedback  <= \s412_feedback ;
    end
    always @(posedge \clk ) begin
        \s414_feedback  <= \s413_feedback ;
    end
    always @(posedge \clk ) begin
        \s415_feedback  <= \s414_feedback ;
    end
    always @(posedge \clk ) begin
        \s416_feedback  <= \s415_feedback ;
    end
    always @(posedge \clk ) begin
        \s417_feedback  <= \s416_feedback ;
    end
    always @(posedge \clk ) begin
        \s418_feedback  <= \s417_feedback ;
    end
    always @(posedge \clk ) begin
        \s419_feedback  <= \s418_feedback ;
    end
    always @(posedge \clk ) begin
        \s420_feedback  <= \s419_feedback ;
    end
    always @(posedge \clk ) begin
        \s421_feedback  <= \s420_feedback ;
    end
    always @(posedge \clk ) begin
        \s422_feedback  <= \s421_feedback ;
    end
    always @(posedge \clk ) begin
        \s423_feedback  <= \s422_feedback ;
    end
    always @(posedge \clk ) begin
        \s424_feedback  <= \s423_feedback ;
    end
    always @(posedge \clk ) begin
        \s425_feedback  <= \s424_feedback ;
    end
    always @(posedge \clk ) begin
        \s426_feedback  <= \s425_feedback ;
    end
    always @(posedge \clk ) begin
        \s427_feedback  <= \s426_feedback ;
    end
    always @(posedge \clk ) begin
        \s428_feedback  <= \s427_feedback ;
    end
    always @(posedge \clk ) begin
        \s429_feedback  <= \s428_feedback ;
    end
    always @(posedge \clk ) begin
        \s430_feedback  <= \s429_feedback ;
    end
    always @(posedge \clk ) begin
        \s431_feedback  <= \s430_feedback ;
    end
    always @(posedge \clk ) begin
        \s432_feedback  <= \s431_feedback ;
    end
    always @(posedge \clk ) begin
        \s433_feedback  <= \s432_feedback ;
    end
    always @(posedge \clk ) begin
        \s434_feedback  <= \s433_feedback ;
    end
    always @(posedge \clk ) begin
        \s435_feedback  <= \s434_feedback ;
    end
    always @(posedge \clk ) begin
        \s436_feedback  <= \s435_feedback ;
    end
    always @(posedge \clk ) begin
        \s437_feedback  <= \s436_feedback ;
    end
    always @(posedge \clk ) begin
        \s438_feedback  <= \s437_feedback ;
    end
    always @(posedge \clk ) begin
        \s439_feedback  <= \s438_feedback ;
    end
    always @(posedge \clk ) begin
        \s440_feedback  <= \s439_feedback ;
    end
    always @(posedge \clk ) begin
        \s441_feedback  <= \s440_feedback ;
    end
    always @(posedge \clk ) begin
        \s442_feedback  <= \s441_feedback ;
    end
    always @(posedge \clk ) begin
        \s443_feedback  <= \s442_feedback ;
    end
    always @(posedge \clk ) begin
        \s444_feedback  <= \s443_feedback ;
    end
    always @(posedge \clk ) begin
        \s445_feedback  <= \s444_feedback ;
    end
    always @(posedge \clk ) begin
        \s446_feedback  <= \s445_feedback ;
    end
    always @(posedge \clk ) begin
        \s447_feedback  <= \s446_feedback ;
    end
    always @(posedge \clk ) begin
        \s448_feedback  <= \s447_feedback ;
    end
    always @(posedge \clk ) begin
        \s449_feedback  <= \s448_feedback ;
    end
    always @(posedge \clk ) begin
        \s450_feedback  <= \s449_feedback ;
    end
    always @(posedge \clk ) begin
        \s451_feedback  <= \s450_feedback ;
    end
    always @(posedge \clk ) begin
        \s452_feedback  <= \s451_feedback ;
    end
    always @(posedge \clk ) begin
        \s453_feedback  <= \s452_feedback ;
    end
    always @(posedge \clk ) begin
        \s454_feedback  <= \s453_feedback ;
    end
    always @(posedge \clk ) begin
        \s455_feedback  <= \s454_feedback ;
    end
    always @(posedge \clk ) begin
        \s456_feedback  <= \s455_feedback ;
    end
    always @(posedge \clk ) begin
        \s457_feedback  <= \s456_feedback ;
    end
    always @(posedge \clk ) begin
        \s458_feedback  <= \s457_feedback ;
    end
    always @(posedge \clk ) begin
        \s459_feedback  <= \s458_feedback ;
    end
    always @(posedge \clk ) begin
        \s460_feedback  <= \s459_feedback ;
    end
    always @(posedge \clk ) begin
        \s461_feedback  <= \s460_feedback ;
    end
    always @(posedge \clk ) begin
        \s462_feedback  <= \s461_feedback ;
    end
    always @(posedge \clk ) begin
        \s463_feedback  <= \s462_feedback ;
    end
    always @(posedge \clk ) begin
        \s464_feedback  <= \s463_feedback ;
    end
    always @(posedge \clk ) begin
        \s465_feedback  <= \s464_feedback ;
    end
    always @(posedge \clk ) begin
        \s466_feedback  <= \s465_feedback ;
    end
    always @(posedge \clk ) begin
        \s467_feedback  <= \s466_feedback ;
    end
    always @(posedge \clk ) begin
        \s468_feedback  <= \s467_feedback ;
    end
    always @(posedge \clk ) begin
        \s469_feedback  <= \s468_feedback ;
    end
    always @(posedge \clk ) begin
        \s470_feedback  <= \s469_feedback ;
    end
    always @(posedge \clk ) begin
        \s471_feedback  <= \s470_feedback ;
    end
    always @(posedge \clk ) begin
        \s472_feedback  <= \s471_feedback ;
    end
    always @(posedge \clk ) begin
        \s473_feedback  <= \s472_feedback ;
    end
    always @(posedge \clk ) begin
        \s474_feedback  <= \s473_feedback ;
    end
    always @(posedge \clk ) begin
        \s475_feedback  <= \s474_feedback ;
    end
    always @(posedge \clk ) begin
        \s476_feedback  <= \s475_feedback ;
    end
    always @(posedge \clk ) begin
        \s477_feedback  <= \s476_feedback ;
    end
    always @(posedge \clk ) begin
        \s478_feedback  <= \s477_feedback ;
    end
    always @(posedge \clk ) begin
        \s479_feedback  <= \s478_feedback ;
    end
    always @(posedge \clk ) begin
        \s480_feedback  <= \s479_feedback ;
    end
    always @(posedge \clk ) begin
        \s481_feedback  <= \s480_feedback ;
    end
    always @(posedge \clk ) begin
        \s482_feedback  <= \s481_feedback ;
    end
    always @(posedge \clk ) begin
        \s483_feedback  <= \s482_feedback ;
    end
    always @(posedge \clk ) begin
        \s484_feedback  <= \s483_feedback ;
    end
    always @(posedge \clk ) begin
        \s485_feedback  <= \s484_feedback ;
    end
    always @(posedge \clk ) begin
        \s486_feedback  <= \s485_feedback ;
    end
    always @(posedge \clk ) begin
        \s487_feedback  <= \s486_feedback ;
    end
    always @(posedge \clk ) begin
        \s488_feedback  <= \s487_feedback ;
    end
    always @(posedge \clk ) begin
        \s489_feedback  <= \s488_feedback ;
    end
    always @(posedge \clk ) begin
        \s490_feedback  <= \s489_feedback ;
    end
    always @(posedge \clk ) begin
        \s491_feedback  <= \s490_feedback ;
    end
    always @(posedge \clk ) begin
        \s492_feedback  <= \s491_feedback ;
    end
    always @(posedge \clk ) begin
        \s493_feedback  <= \s492_feedback ;
    end
    always @(posedge \clk ) begin
        \s494_feedback  <= \s493_feedback ;
    end
    always @(posedge \clk ) begin
        \s495_feedback  <= \s494_feedback ;
    end
    always @(posedge \clk ) begin
        \s496_feedback  <= \s495_feedback ;
    end
    always @(posedge \clk ) begin
        \s497_feedback  <= \s496_feedback ;
    end
    always @(posedge \clk ) begin
        \s498_feedback  <= \s497_feedback ;
    end
    always @(posedge \clk ) begin
        \s499_feedback  <= \s498_feedback ;
    end
    always @(posedge \clk ) begin
        \s500_feedback  <= \s499_feedback ;
    end
    always @(posedge \clk ) begin
        \s501_feedback  <= \s500_feedback ;
    end
    always @(posedge \clk ) begin
        \s502_feedback  <= \s501_feedback ;
    end
    always @(posedge \clk ) begin
        \s503_feedback  <= \s502_feedback ;
    end
    always @(posedge \clk ) begin
        \s504_feedback  <= \s503_feedback ;
    end
    always @(posedge \clk ) begin
        \s505_feedback  <= \s504_feedback ;
    end
    always @(posedge \clk ) begin
        \s506_feedback  <= \s505_feedback ;
    end
    always @(posedge \clk ) begin
        \s507_feedback  <= \s506_feedback ;
    end
    always @(posedge \clk ) begin
        \s508_feedback  <= \s507_feedback ;
    end
    always @(posedge \clk ) begin
        \s509_feedback  <= \s508_feedback ;
    end
    always @(posedge \clk ) begin
        \s510_feedback  <= \s509_feedback ;
    end
    always @(posedge \clk ) begin
        \s511_feedback  <= \s510_feedback ;
    end
    always @(posedge \clk ) begin
        \s512_feedback  <= \s511_feedback ;
    end
    always @(posedge \clk ) begin
        \s513_feedback  <= \s512_feedback ;
    end
    always @(posedge \clk ) begin
        \s514_feedback  <= \s513_feedback ;
    end
    always @(posedge \clk ) begin
        \s515_feedback  <= \s514_feedback ;
    end
    always @(posedge \clk ) begin
        \s516_feedback  <= \s515_feedback ;
    end
    always @(posedge \clk ) begin
        \s517_feedback  <= \s516_feedback ;
    end
    always @(posedge \clk ) begin
        \s518_feedback  <= \s517_feedback ;
    end
    always @(posedge \clk ) begin
        \s519_feedback  <= \s518_feedback ;
    end
    always @(posedge \clk ) begin
        \s520_feedback  <= \s519_feedback ;
    end
    always @(posedge \clk ) begin
        \s521_feedback  <= \s520_feedback ;
    end
    always @(posedge \clk ) begin
        \s522_feedback  <= \s521_feedback ;
    end
    always @(posedge \clk ) begin
        \s523_feedback  <= \s522_feedback ;
    end
    always @(posedge \clk ) begin
        \s524_feedback  <= \s523_feedback ;
    end
    always @(posedge \clk ) begin
        \s525_feedback  <= \s524_feedback ;
    end
    always @(posedge \clk ) begin
        \s526_feedback  <= \s525_feedback ;
    end
    always @(posedge \clk ) begin
        \s527_feedback  <= \s526_feedback ;
    end
    always @(posedge \clk ) begin
        \s528_feedback  <= \s527_feedback ;
    end
    always @(posedge \clk ) begin
        \s529_feedback  <= \s528_feedback ;
    end
    always @(posedge \clk ) begin
        \s530_feedback  <= \s529_feedback ;
    end
    always @(posedge \clk ) begin
        \s531_feedback  <= \s530_feedback ;
    end
    always @(posedge \clk ) begin
        \s532_feedback  <= \s531_feedback ;
    end
    always @(posedge \clk ) begin
        \s533_feedback  <= \s532_feedback ;
    end
    always @(posedge \clk ) begin
        \s534_feedback  <= \s533_feedback ;
    end
    always @(posedge \clk ) begin
        \s535_feedback  <= \s534_feedback ;
    end
    always @(posedge \clk ) begin
        \s536_feedback  <= \s535_feedback ;
    end
    always @(posedge \clk ) begin
        \s537_feedback  <= \s536_feedback ;
    end
    always @(posedge \clk ) begin
        \s538_feedback  <= \s537_feedback ;
    end
    always @(posedge \clk ) begin
        \s539_feedback  <= \s538_feedback ;
    end
    always @(posedge \clk ) begin
        \s540_feedback  <= \s539_feedback ;
    end
    always @(posedge \clk ) begin
        \s541_feedback  <= \s540_feedback ;
    end
    always @(posedge \clk ) begin
        \s542_feedback  <= \s541_feedback ;
    end
    always @(posedge \clk ) begin
        \s543_feedback  <= \s542_feedback ;
    end
    always @(posedge \clk ) begin
        \s544_feedback  <= \s543_feedback ;
    end
    always @(posedge \clk ) begin
        \s545_feedback  <= \s544_feedback ;
    end
    always @(posedge \clk ) begin
        \s546_feedback  <= \s545_feedback ;
    end
    always @(posedge \clk ) begin
        \s547_feedback  <= \s546_feedback ;
    end
    always @(posedge \clk ) begin
        \s548_feedback  <= \s547_feedback ;
    end
    always @(posedge \clk ) begin
        \s549_feedback  <= \s548_feedback ;
    end
    always @(posedge \clk ) begin
        \s550_feedback  <= \s549_feedback ;
    end
    always @(posedge \clk ) begin
        \s551_feedback  <= \s550_feedback ;
    end
    always @(posedge \clk ) begin
        \s552_feedback  <= \s551_feedback ;
    end
    always @(posedge \clk ) begin
        \s553_feedback  <= \s552_feedback ;
    end
    always @(posedge \clk ) begin
        \s554_feedback  <= \s553_feedback ;
    end
    always @(posedge \clk ) begin
        \s555_feedback  <= \s554_feedback ;
    end
    always @(posedge \clk ) begin
        \s556_feedback  <= \s555_feedback ;
    end
    always @(posedge \clk ) begin
        \s557_feedback  <= \s556_feedback ;
    end
    always @(posedge \clk ) begin
        \s558_feedback  <= \s557_feedback ;
    end
    always @(posedge \clk ) begin
        \s559_feedback  <= \s558_feedback ;
    end
    always @(posedge \clk ) begin
        \s560_feedback  <= \s559_feedback ;
    end
    always @(posedge \clk ) begin
        \s561_feedback  <= \s560_feedback ;
    end
    always @(posedge \clk ) begin
        \s562_feedback  <= \s561_feedback ;
    end
    always @(posedge \clk ) begin
        \s563_feedback  <= \s562_feedback ;
    end
    always @(posedge \clk ) begin
        \s564_feedback  <= \s563_feedback ;
    end
    always @(posedge \clk ) begin
        \s565_feedback  <= \s564_feedback ;
    end
    always @(posedge \clk ) begin
        \s566_feedback  <= \s565_feedback ;
    end
    always @(posedge \clk ) begin
        \s567_feedback  <= \s566_feedback ;
    end
    always @(posedge \clk ) begin
        \s568_feedback  <= \s567_feedback ;
    end
    always @(posedge \clk ) begin
        \s569_feedback  <= \s568_feedback ;
    end
    always @(posedge \clk ) begin
        \s570_feedback  <= \s569_feedback ;
    end
    always @(posedge \clk ) begin
        \s571_feedback  <= \s570_feedback ;
    end
    always @(posedge \clk ) begin
        \s572_feedback  <= \s571_feedback ;
    end
    always @(posedge \clk ) begin
        \s573_feedback  <= \s572_feedback ;
    end
    always @(posedge \clk ) begin
        \s574_feedback  <= \s573_feedback ;
    end
    always @(posedge \clk ) begin
        \s575_feedback  <= \s574_feedback ;
    end
    always @(posedge \clk ) begin
        \s576_feedback  <= \s575_feedback ;
    end
    always @(posedge \clk ) begin
        \s577_feedback  <= \s576_feedback ;
    end
    always @(posedge \clk ) begin
        \s578_feedback  <= \s577_feedback ;
    end
    always @(posedge \clk ) begin
        \s579_feedback  <= \s578_feedback ;
    end
    always @(posedge \clk ) begin
        \s580_feedback  <= \s579_feedback ;
    end
    always @(posedge \clk ) begin
        \s581_feedback  <= \s580_feedback ;
    end
    always @(posedge \clk ) begin
        \s582_feedback  <= \s581_feedback ;
    end
    always @(posedge \clk ) begin
        \s583_feedback  <= \s582_feedback ;
    end
    always @(posedge \clk ) begin
        \s584_feedback  <= \s583_feedback ;
    end
    always @(posedge \clk ) begin
        \s585_feedback  <= \s584_feedback ;
    end
    always @(posedge \clk ) begin
        \s586_feedback  <= \s585_feedback ;
    end
    always @(posedge \clk ) begin
        \s587_feedback  <= \s586_feedback ;
    end
    always @(posedge \clk ) begin
        \s588_feedback  <= \s587_feedback ;
    end
    always @(posedge \clk ) begin
        \s589_feedback  <= \s588_feedback ;
    end
    always @(posedge \clk ) begin
        \s590_feedback  <= \s589_feedback ;
    end
    always @(posedge \clk ) begin
        \s591_feedback  <= \s590_feedback ;
    end
    always @(posedge \clk ) begin
        \s592_feedback  <= \s591_feedback ;
    end
    always @(posedge \clk ) begin
        \s593_feedback  <= \s592_feedback ;
    end
    always @(posedge \clk ) begin
        \s594_feedback  <= \s593_feedback ;
    end
    always @(posedge \clk ) begin
        \s595_feedback  <= \s594_feedback ;
    end
    always @(posedge \clk ) begin
        \s596_feedback  <= \s595_feedback ;
    end
    always @(posedge \clk ) begin
        \s597_feedback  <= \s596_feedback ;
    end
    always @(posedge \clk ) begin
        \s598_feedback  <= \s597_feedback ;
    end
    always @(posedge \clk ) begin
        \s599_feedback  <= \s598_feedback ;
    end
    always @(posedge \clk ) begin
        \s600_feedback  <= \s599_feedback ;
    end
    assign output__ = \s600_feedback ;
endmodule

module tt_um_delay_line_tmng (
        input[7:0] ui_in,
        output[7:0] uo_out,
        input[7:0] uio_in,
        output[7:0] uio_out,
        output[7:0] uio_oe,
        input ena,
        input clk,
        input rst_n
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "tt_um_delay_line_tmng" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, tt_um_delay_line_tmng);
        end
    end
    `endif
    logic[7:0] \uo_out_mut ;
    assign uo_out = \uo_out_mut ;
    logic[7:0] \uio_out_mut ;
    assign uio_out = \uio_out_mut ;
    logic[7:0] \uio_oe_mut ;
    assign uio_oe = \uio_oe_mut ;
    (* src = "src/main.spade:25,38" *)
    logic[7:0] _e_623;
    logic[2:0] _e_625;
    (* src = "src/main.spade:25,38" *)
    logic _e_622;
    (* src = "src/main.spade:25,13" *)
    logic \x ;
    logic[7:0] _e_631;
    logic[7:0] _e_633;
    (* src = "src/main.spade:28,18" *)
    logic[7:0] _e_628;
    logic[7:0] _e_635;
    logic[7:0] _e_637;
    (* src = "src/main.spade:25,38" *)
    \std::conv::int_to_bits[1546]  int_to_bits_0(.input_i(\ui_in ), .output__(_e_623));
    assign _e_625 = 0;
    assign _e_622 = _e_623[_e_625];
    (* src = "src/main.spade:25,13" *)
    \tt07_delay_line_tmng::main::shift_reg  shift_reg_0(.clk_i(\clk ), .feedback_i(_e_622), .output__(\x ));
    assign _e_631 = 1;
    assign _e_633 = 0;
    assign _e_628 = \x  ? _e_631 : _e_633;
    assign \uo_out_mut  = _e_628;
    assign _e_635 = 0;
    assign \uio_out_mut  = _e_635;
    assign _e_637 = 0;
    assign \uio_oe_mut  = _e_637;
endmodule

module \std::cdc::unsafe::sync2[345]  (
        input clk_i,
        input in_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::cdc::unsafe::sync2[345]" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::cdc::unsafe::sync2[345] );
        end
    end
    `endif
    logic \clk ;
    assign \clk  = clk_i;
    logic \in ;
    assign \in  = in_i;
    (* src = "<compiler dir>/stdlib/cdc.spade:20,18" *)
    reg \sync1 ;
    (* src = "<compiler dir>/stdlib/cdc.spade:21,18" *)
    reg \sync2 ;
    always @(posedge \clk ) begin
        \sync1  <= \in ;
    end
    always @(posedge \clk ) begin
        \sync2  <= \sync1 ;
    end
    assign output__ = \sync2 ;
endmodule

module \std::conv::int_to_bits[1546]  (
        input[7:0] input_i,
        output[7:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::int_to_bits[1546]" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::int_to_bits[1546] );
        end
    end
    `endif
    logic[7:0] \input ;
    assign \input  = input_i;
    logic[7:0] _e_4;
    assign _e_4 = \input ;
    assign output__ = _e_4;
endmodule