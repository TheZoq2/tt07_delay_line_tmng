module \std::conv::bit_to_bool  (
        input b_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::bit_to_bool" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::bit_to_bool );
        end
    end
    `endif
    logic \b ;
    assign \b  = b_i;
    logic _e_1;
    assign _e_1 = \b ;
    assign output__ = _e_1;
endmodule

module \std::conv::unsafe::clock_to_bool  (
        input c_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::unsafe::clock_to_bool" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::unsafe::clock_to_bool );
        end
    end
    `endif
    logic \c ;
    assign \c  = c_i;
    logic _e_22;
    assign _e_22 = \c ;
    assign output__ = _e_22;
endmodule

module \std::conv::unsafe::bool_to_clock  (
        input c_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::unsafe::bool_to_clock" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::unsafe::bool_to_clock );
        end
    end
    `endif
    logic \c ;
    assign \c  = c_i;
    logic _e_25;
    assign _e_25 = \c ;
    assign output__ = _e_25;
endmodule

module \std::io::rising_edge  (
        input clk_i,
        input sync1_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::io::rising_edge" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::io::rising_edge );
        end
    end
    `endif
    logic \clk ;
    assign \clk  = clk_i;
    logic \sync1 ;
    assign \sync1  = sync1_i;
    (* src = "<compiler dir>/stdlib/io.spade:3,14" *)
    reg \sync2 ;
    (* src = "<compiler dir>/stdlib/io.spade:4,14" *)
    logic _e_33;
    (* src = "<compiler dir>/stdlib/io.spade:4,5" *)
    logic _e_31;
    always @(posedge \clk ) begin
        \sync2  <= \sync1 ;
    end
    assign _e_33 = !\sync2 ;
    assign _e_31 = \sync1  && _e_33;
    assign output__ = _e_31;
endmodule

module \std::io::falling_edge  (
        input clk_i,
        input sync1_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::io::falling_edge" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::io::falling_edge );
        end
    end
    `endif
    logic \clk ;
    assign \clk  = clk_i;
    logic \sync1 ;
    assign \sync1  = sync1_i;
    (* src = "<compiler dir>/stdlib/io.spade:9,14" *)
    reg \sync2 ;
    (* src = "<compiler dir>/stdlib/io.spade:10,14" *)
    logic _e_41;
    (* src = "<compiler dir>/stdlib/io.spade:10,5" *)
    logic _e_39;
    always @(posedge \clk ) begin
        \sync2  <= \sync1 ;
    end
    assign _e_41 = !\sync1 ;
    assign _e_39 = \sync2  && _e_41;
    assign output__ = _e_39;
endmodule

module \std::cdc::sync2_bool  (
        input clk_i,
        input in_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::cdc::sync2_bool" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::cdc::sync2_bool );
        end
    end
    `endif
    logic \clk ;
    assign \clk  = clk_i;
    logic \in ;
    assign \in  = in_i;
    (* src = "<compiler dir>/stdlib/cdc.spade:38,5" *)
    logic _e_335;
    (* src = "<compiler dir>/stdlib/cdc.spade:38,5" *)
    \std::cdc::unsafe::sync2[431]  sync2_0(.clk_i(\clk ), .in_i(\in ), .output__(_e_335));
    assign output__ = _e_335;
endmodule

module \tt07_delay_line_tmng::sreg::dlygate  (
        input A_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "tt07_delay_line_tmng::sreg::dlygate" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \tt07_delay_line_tmng::sreg::dlygate );
        end
    end
    `endif
    logic \A ;
    assign \A  = A_i;
    logic \X_mut ;
    logic _e_624;
    
    (* src = "src/sreg.spade:9,13" *)
    sky130_fd_sc_hd__dlygate4sd1_1 sky130_fd_sc_hd__dlygate4sd1_1_0(.A(\A ), .X(\X_mut ));
    assign _e_624 = \X_mut ;
    assign output__ = _e_624;
endmodule

module \tt07_delay_line_tmng::sreg::inv_reg  (
        input clk_i,
        input val_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "tt07_delay_line_tmng::sreg::inv_reg" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \tt07_delay_line_tmng::sreg::inv_reg );
        end
    end
    `endif
    logic \clk ;
    assign \clk  = clk_i;
    logic \val ;
    assign \val  = val_i;
    (* src = "src/sreg.spade:16,5" *)
    reg \s1_val ;
    (* src = "src/sreg.spade:16,5" *)
    reg s1_val_n1;
    (* src = "src/sreg.spade:18,5" *)
    reg \s2_val ;
    (* src = "src/sreg.spade:18,5" *)
    reg s2_val_n1;
    (* src = "src/sreg.spade:18,5" *)
    reg s2_val_n2;
    (* src = "src/sreg.spade:15,19" *)
    logic val_n1;
    (* src = "src/sreg.spade:17,19" *)
    logic val_n2;
    always @(posedge \clk ) begin
        \s1_val  <= \val ;
    end
    always @(posedge \clk ) begin
        s1_val_n1 <= val_n1;
    end
    always @(posedge \clk ) begin
        \s2_val  <= \s1_val ;
    end
    always @(posedge \clk ) begin
        s2_val_n1 <= s1_val_n1;
    end
    always @(posedge \clk ) begin
        s2_val_n2 <= val_n2;
    end
    (* src = "src/sreg.spade:15,19" *)
    \tt07_delay_line_tmng::sreg::dlygate  dlygate_0(.A_i(\val ), .output__(val_n1));
    (* src = "src/sreg.spade:17,19" *)
    \tt07_delay_line_tmng::sreg::dlygate  dlygate_1(.A_i(s1_val_n1), .output__(val_n2));
    assign output__ = s2_val_n2;
endmodule

module \tt07_delay_line_tmng::sreg::shift_reg100  (
        input clk_i,
        input val_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "tt07_delay_line_tmng::sreg::shift_reg100" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \tt07_delay_line_tmng::sreg::shift_reg100 );
        end
    end
    `endif
    logic \clk ;
    assign \clk  = clk_i;
    logic \val ;
    assign \val  = val_i;
    (* src = "src/sreg.spade:24,5" *)
    reg \s1_val ;
    (* src = "src/sreg.spade:24,5" *)
    reg \s2_val ;
    (* src = "src/sreg.spade:26,5" *)
    reg \s3_val ;
    (* src = "src/sreg.spade:26,5" *)
    reg \s4_val ;
    (* src = "src/sreg.spade:28,5" *)
    reg \s5_val ;
    (* src = "src/sreg.spade:28,5" *)
    reg s5_val_n1;
    (* src = "src/sreg.spade:28,5" *)
    reg \s6_val ;
    (* src = "src/sreg.spade:28,5" *)
    reg s6_val_n1;
    (* src = "src/sreg.spade:30,5" *)
    reg \s7_val ;
    (* src = "src/sreg.spade:30,5" *)
    reg s7_val_n1;
    (* src = "src/sreg.spade:30,5" *)
    reg s7_val_n2;
    (* src = "src/sreg.spade:30,5" *)
    reg \s8_val ;
    (* src = "src/sreg.spade:30,5" *)
    reg s8_val_n1;
    (* src = "src/sreg.spade:30,5" *)
    reg s8_val_n2;
    (* src = "src/sreg.spade:32,5" *)
    reg \s9_val ;
    (* src = "src/sreg.spade:32,5" *)
    reg s9_val_n1;
    (* src = "src/sreg.spade:32,5" *)
    reg s9_val_n2;
    (* src = "src/sreg.spade:32,5" *)
    reg s9_val_n3;
    (* src = "src/sreg.spade:32,5" *)
    reg \s10_val ;
    (* src = "src/sreg.spade:32,5" *)
    reg s10_val_n1;
    (* src = "src/sreg.spade:32,5" *)
    reg s10_val_n2;
    (* src = "src/sreg.spade:32,5" *)
    reg s10_val_n3;
    (* src = "src/sreg.spade:34,5" *)
    reg \s11_val ;
    (* src = "src/sreg.spade:34,5" *)
    reg s11_val_n1;
    (* src = "src/sreg.spade:34,5" *)
    reg s11_val_n2;
    (* src = "src/sreg.spade:34,5" *)
    reg s11_val_n3;
    (* src = "src/sreg.spade:34,5" *)
    reg s11_val_n4;
    (* src = "src/sreg.spade:34,5" *)
    reg \s12_val ;
    (* src = "src/sreg.spade:34,5" *)
    reg s12_val_n1;
    (* src = "src/sreg.spade:34,5" *)
    reg s12_val_n2;
    (* src = "src/sreg.spade:34,5" *)
    reg s12_val_n3;
    (* src = "src/sreg.spade:34,5" *)
    reg s12_val_n4;
    (* src = "src/sreg.spade:36,5" *)
    reg \s13_val ;
    (* src = "src/sreg.spade:36,5" *)
    reg s13_val_n1;
    (* src = "src/sreg.spade:36,5" *)
    reg s13_val_n2;
    (* src = "src/sreg.spade:36,5" *)
    reg s13_val_n3;
    (* src = "src/sreg.spade:36,5" *)
    reg s13_val_n4;
    (* src = "src/sreg.spade:36,5" *)
    reg s13_val_n5;
    (* src = "src/sreg.spade:36,5" *)
    reg \s14_val ;
    (* src = "src/sreg.spade:36,5" *)
    reg s14_val_n1;
    (* src = "src/sreg.spade:36,5" *)
    reg s14_val_n2;
    (* src = "src/sreg.spade:36,5" *)
    reg s14_val_n3;
    (* src = "src/sreg.spade:36,5" *)
    reg s14_val_n4;
    (* src = "src/sreg.spade:36,5" *)
    reg s14_val_n5;
    (* src = "src/sreg.spade:38,5" *)
    reg \s15_val ;
    (* src = "src/sreg.spade:38,5" *)
    reg s15_val_n1;
    (* src = "src/sreg.spade:38,5" *)
    reg s15_val_n2;
    (* src = "src/sreg.spade:38,5" *)
    reg s15_val_n3;
    (* src = "src/sreg.spade:38,5" *)
    reg s15_val_n4;
    (* src = "src/sreg.spade:38,5" *)
    reg s15_val_n5;
    (* src = "src/sreg.spade:38,5" *)
    reg s15_val_n6;
    (* src = "src/sreg.spade:38,5" *)
    reg \s16_val ;
    (* src = "src/sreg.spade:38,5" *)
    reg s16_val_n1;
    (* src = "src/sreg.spade:38,5" *)
    reg s16_val_n2;
    (* src = "src/sreg.spade:38,5" *)
    reg s16_val_n3;
    (* src = "src/sreg.spade:38,5" *)
    reg s16_val_n4;
    (* src = "src/sreg.spade:38,5" *)
    reg s16_val_n5;
    (* src = "src/sreg.spade:38,5" *)
    reg s16_val_n6;
    (* src = "src/sreg.spade:40,5" *)
    reg \s17_val ;
    (* src = "src/sreg.spade:40,5" *)
    reg s17_val_n1;
    (* src = "src/sreg.spade:40,5" *)
    reg s17_val_n2;
    (* src = "src/sreg.spade:40,5" *)
    reg s17_val_n3;
    (* src = "src/sreg.spade:40,5" *)
    reg s17_val_n4;
    (* src = "src/sreg.spade:40,5" *)
    reg s17_val_n5;
    (* src = "src/sreg.spade:40,5" *)
    reg s17_val_n6;
    (* src = "src/sreg.spade:40,5" *)
    reg s17_val_n7;
    (* src = "src/sreg.spade:40,5" *)
    reg \s18_val ;
    (* src = "src/sreg.spade:40,5" *)
    reg s18_val_n1;
    (* src = "src/sreg.spade:40,5" *)
    reg s18_val_n2;
    (* src = "src/sreg.spade:40,5" *)
    reg s18_val_n3;
    (* src = "src/sreg.spade:40,5" *)
    reg s18_val_n4;
    (* src = "src/sreg.spade:40,5" *)
    reg s18_val_n5;
    (* src = "src/sreg.spade:40,5" *)
    reg s18_val_n6;
    (* src = "src/sreg.spade:40,5" *)
    reg s18_val_n7;
    (* src = "src/sreg.spade:42,5" *)
    reg \s19_val ;
    (* src = "src/sreg.spade:42,5" *)
    reg s19_val_n1;
    (* src = "src/sreg.spade:42,5" *)
    reg s19_val_n2;
    (* src = "src/sreg.spade:42,5" *)
    reg s19_val_n3;
    (* src = "src/sreg.spade:42,5" *)
    reg s19_val_n4;
    (* src = "src/sreg.spade:42,5" *)
    reg s19_val_n5;
    (* src = "src/sreg.spade:42,5" *)
    reg s19_val_n6;
    (* src = "src/sreg.spade:42,5" *)
    reg s19_val_n7;
    (* src = "src/sreg.spade:42,5" *)
    reg s19_val_n8;
    (* src = "src/sreg.spade:42,5" *)
    reg \s20_val ;
    (* src = "src/sreg.spade:42,5" *)
    reg s20_val_n1;
    (* src = "src/sreg.spade:42,5" *)
    reg s20_val_n2;
    (* src = "src/sreg.spade:42,5" *)
    reg s20_val_n3;
    (* src = "src/sreg.spade:42,5" *)
    reg s20_val_n4;
    (* src = "src/sreg.spade:42,5" *)
    reg s20_val_n5;
    (* src = "src/sreg.spade:42,5" *)
    reg s20_val_n6;
    (* src = "src/sreg.spade:42,5" *)
    reg s20_val_n7;
    (* src = "src/sreg.spade:42,5" *)
    reg s20_val_n8;
    (* src = "src/sreg.spade:44,5" *)
    reg \s21_val ;
    (* src = "src/sreg.spade:44,5" *)
    reg s21_val_n1;
    (* src = "src/sreg.spade:44,5" *)
    reg s21_val_n2;
    (* src = "src/sreg.spade:44,5" *)
    reg s21_val_n3;
    (* src = "src/sreg.spade:44,5" *)
    reg s21_val_n4;
    (* src = "src/sreg.spade:44,5" *)
    reg s21_val_n5;
    (* src = "src/sreg.spade:44,5" *)
    reg s21_val_n6;
    (* src = "src/sreg.spade:44,5" *)
    reg s21_val_n7;
    (* src = "src/sreg.spade:44,5" *)
    reg s21_val_n8;
    (* src = "src/sreg.spade:44,5" *)
    reg s21_val_n9;
    (* src = "src/sreg.spade:44,5" *)
    reg \s22_val ;
    (* src = "src/sreg.spade:44,5" *)
    reg s22_val_n1;
    (* src = "src/sreg.spade:44,5" *)
    reg s22_val_n2;
    (* src = "src/sreg.spade:44,5" *)
    reg s22_val_n3;
    (* src = "src/sreg.spade:44,5" *)
    reg s22_val_n4;
    (* src = "src/sreg.spade:44,5" *)
    reg s22_val_n5;
    (* src = "src/sreg.spade:44,5" *)
    reg s22_val_n6;
    (* src = "src/sreg.spade:44,5" *)
    reg s22_val_n7;
    (* src = "src/sreg.spade:44,5" *)
    reg s22_val_n8;
    (* src = "src/sreg.spade:44,5" *)
    reg s22_val_n9;
    (* src = "src/sreg.spade:46,5" *)
    reg \s23_val ;
    (* src = "src/sreg.spade:46,5" *)
    reg s23_val_n1;
    (* src = "src/sreg.spade:46,5" *)
    reg s23_val_n2;
    (* src = "src/sreg.spade:46,5" *)
    reg s23_val_n3;
    (* src = "src/sreg.spade:46,5" *)
    reg s23_val_n4;
    (* src = "src/sreg.spade:46,5" *)
    reg s23_val_n5;
    (* src = "src/sreg.spade:46,5" *)
    reg s23_val_n6;
    (* src = "src/sreg.spade:46,5" *)
    reg s23_val_n7;
    (* src = "src/sreg.spade:46,5" *)
    reg s23_val_n8;
    (* src = "src/sreg.spade:46,5" *)
    reg s23_val_n9;
    (* src = "src/sreg.spade:46,5" *)
    reg s23_val_n10;
    (* src = "src/sreg.spade:46,5" *)
    reg \s24_val ;
    (* src = "src/sreg.spade:46,5" *)
    reg s24_val_n1;
    (* src = "src/sreg.spade:46,5" *)
    reg s24_val_n2;
    (* src = "src/sreg.spade:46,5" *)
    reg s24_val_n3;
    (* src = "src/sreg.spade:46,5" *)
    reg s24_val_n4;
    (* src = "src/sreg.spade:46,5" *)
    reg s24_val_n5;
    (* src = "src/sreg.spade:46,5" *)
    reg s24_val_n6;
    (* src = "src/sreg.spade:46,5" *)
    reg s24_val_n7;
    (* src = "src/sreg.spade:46,5" *)
    reg s24_val_n8;
    (* src = "src/sreg.spade:46,5" *)
    reg s24_val_n9;
    (* src = "src/sreg.spade:46,5" *)
    reg s24_val_n10;
    (* src = "src/sreg.spade:48,5" *)
    reg \s25_val ;
    (* src = "src/sreg.spade:48,5" *)
    reg s25_val_n1;
    (* src = "src/sreg.spade:48,5" *)
    reg s25_val_n2;
    (* src = "src/sreg.spade:48,5" *)
    reg s25_val_n3;
    (* src = "src/sreg.spade:48,5" *)
    reg s25_val_n4;
    (* src = "src/sreg.spade:48,5" *)
    reg s25_val_n5;
    (* src = "src/sreg.spade:48,5" *)
    reg s25_val_n6;
    (* src = "src/sreg.spade:48,5" *)
    reg s25_val_n7;
    (* src = "src/sreg.spade:48,5" *)
    reg s25_val_n8;
    (* src = "src/sreg.spade:48,5" *)
    reg s25_val_n9;
    (* src = "src/sreg.spade:48,5" *)
    reg s25_val_n10;
    (* src = "src/sreg.spade:48,5" *)
    reg s25_val_n11;
    (* src = "src/sreg.spade:48,5" *)
    reg \s26_val ;
    (* src = "src/sreg.spade:48,5" *)
    reg s26_val_n1;
    (* src = "src/sreg.spade:48,5" *)
    reg s26_val_n2;
    (* src = "src/sreg.spade:48,5" *)
    reg s26_val_n3;
    (* src = "src/sreg.spade:48,5" *)
    reg s26_val_n4;
    (* src = "src/sreg.spade:48,5" *)
    reg s26_val_n5;
    (* src = "src/sreg.spade:48,5" *)
    reg s26_val_n6;
    (* src = "src/sreg.spade:48,5" *)
    reg s26_val_n7;
    (* src = "src/sreg.spade:48,5" *)
    reg s26_val_n8;
    (* src = "src/sreg.spade:48,5" *)
    reg s26_val_n9;
    (* src = "src/sreg.spade:48,5" *)
    reg s26_val_n10;
    (* src = "src/sreg.spade:48,5" *)
    reg s26_val_n11;
    (* src = "src/sreg.spade:50,5" *)
    reg \s27_val ;
    (* src = "src/sreg.spade:50,5" *)
    reg s27_val_n1;
    (* src = "src/sreg.spade:50,5" *)
    reg s27_val_n2;
    (* src = "src/sreg.spade:50,5" *)
    reg s27_val_n3;
    (* src = "src/sreg.spade:50,5" *)
    reg s27_val_n4;
    (* src = "src/sreg.spade:50,5" *)
    reg s27_val_n5;
    (* src = "src/sreg.spade:50,5" *)
    reg s27_val_n6;
    (* src = "src/sreg.spade:50,5" *)
    reg s27_val_n7;
    (* src = "src/sreg.spade:50,5" *)
    reg s27_val_n8;
    (* src = "src/sreg.spade:50,5" *)
    reg s27_val_n9;
    (* src = "src/sreg.spade:50,5" *)
    reg s27_val_n10;
    (* src = "src/sreg.spade:50,5" *)
    reg s27_val_n11;
    (* src = "src/sreg.spade:50,5" *)
    reg s27_val_n12;
    (* src = "src/sreg.spade:50,5" *)
    reg \s28_val ;
    (* src = "src/sreg.spade:50,5" *)
    reg s28_val_n1;
    (* src = "src/sreg.spade:50,5" *)
    reg s28_val_n2;
    (* src = "src/sreg.spade:50,5" *)
    reg s28_val_n3;
    (* src = "src/sreg.spade:50,5" *)
    reg s28_val_n4;
    (* src = "src/sreg.spade:50,5" *)
    reg s28_val_n5;
    (* src = "src/sreg.spade:50,5" *)
    reg s28_val_n6;
    (* src = "src/sreg.spade:50,5" *)
    reg s28_val_n7;
    (* src = "src/sreg.spade:50,5" *)
    reg s28_val_n8;
    (* src = "src/sreg.spade:50,5" *)
    reg s28_val_n9;
    (* src = "src/sreg.spade:50,5" *)
    reg s28_val_n10;
    (* src = "src/sreg.spade:50,5" *)
    reg s28_val_n11;
    (* src = "src/sreg.spade:50,5" *)
    reg s28_val_n12;
    (* src = "src/sreg.spade:52,5" *)
    reg \s29_val ;
    (* src = "src/sreg.spade:52,5" *)
    reg s29_val_n1;
    (* src = "src/sreg.spade:52,5" *)
    reg s29_val_n2;
    (* src = "src/sreg.spade:52,5" *)
    reg s29_val_n3;
    (* src = "src/sreg.spade:52,5" *)
    reg s29_val_n4;
    (* src = "src/sreg.spade:52,5" *)
    reg s29_val_n5;
    (* src = "src/sreg.spade:52,5" *)
    reg s29_val_n6;
    (* src = "src/sreg.spade:52,5" *)
    reg s29_val_n7;
    (* src = "src/sreg.spade:52,5" *)
    reg s29_val_n8;
    (* src = "src/sreg.spade:52,5" *)
    reg s29_val_n9;
    (* src = "src/sreg.spade:52,5" *)
    reg s29_val_n10;
    (* src = "src/sreg.spade:52,5" *)
    reg s29_val_n11;
    (* src = "src/sreg.spade:52,5" *)
    reg s29_val_n12;
    (* src = "src/sreg.spade:52,5" *)
    reg s29_val_n13;
    (* src = "src/sreg.spade:52,5" *)
    reg \s30_val ;
    (* src = "src/sreg.spade:52,5" *)
    reg s30_val_n1;
    (* src = "src/sreg.spade:52,5" *)
    reg s30_val_n2;
    (* src = "src/sreg.spade:52,5" *)
    reg s30_val_n3;
    (* src = "src/sreg.spade:52,5" *)
    reg s30_val_n4;
    (* src = "src/sreg.spade:52,5" *)
    reg s30_val_n5;
    (* src = "src/sreg.spade:52,5" *)
    reg s30_val_n6;
    (* src = "src/sreg.spade:52,5" *)
    reg s30_val_n7;
    (* src = "src/sreg.spade:52,5" *)
    reg s30_val_n8;
    (* src = "src/sreg.spade:52,5" *)
    reg s30_val_n9;
    (* src = "src/sreg.spade:52,5" *)
    reg s30_val_n10;
    (* src = "src/sreg.spade:52,5" *)
    reg s30_val_n11;
    (* src = "src/sreg.spade:52,5" *)
    reg s30_val_n12;
    (* src = "src/sreg.spade:52,5" *)
    reg s30_val_n13;
    (* src = "src/sreg.spade:54,5" *)
    reg \s31_val ;
    (* src = "src/sreg.spade:54,5" *)
    reg s31_val_n1;
    (* src = "src/sreg.spade:54,5" *)
    reg s31_val_n2;
    (* src = "src/sreg.spade:54,5" *)
    reg s31_val_n3;
    (* src = "src/sreg.spade:54,5" *)
    reg s31_val_n4;
    (* src = "src/sreg.spade:54,5" *)
    reg s31_val_n5;
    (* src = "src/sreg.spade:54,5" *)
    reg s31_val_n6;
    (* src = "src/sreg.spade:54,5" *)
    reg s31_val_n7;
    (* src = "src/sreg.spade:54,5" *)
    reg s31_val_n8;
    (* src = "src/sreg.spade:54,5" *)
    reg s31_val_n9;
    (* src = "src/sreg.spade:54,5" *)
    reg s31_val_n10;
    (* src = "src/sreg.spade:54,5" *)
    reg s31_val_n11;
    (* src = "src/sreg.spade:54,5" *)
    reg s31_val_n12;
    (* src = "src/sreg.spade:54,5" *)
    reg s31_val_n13;
    (* src = "src/sreg.spade:54,5" *)
    reg s31_val_n14;
    (* src = "src/sreg.spade:54,5" *)
    reg \s32_val ;
    (* src = "src/sreg.spade:54,5" *)
    reg s32_val_n1;
    (* src = "src/sreg.spade:54,5" *)
    reg s32_val_n2;
    (* src = "src/sreg.spade:54,5" *)
    reg s32_val_n3;
    (* src = "src/sreg.spade:54,5" *)
    reg s32_val_n4;
    (* src = "src/sreg.spade:54,5" *)
    reg s32_val_n5;
    (* src = "src/sreg.spade:54,5" *)
    reg s32_val_n6;
    (* src = "src/sreg.spade:54,5" *)
    reg s32_val_n7;
    (* src = "src/sreg.spade:54,5" *)
    reg s32_val_n8;
    (* src = "src/sreg.spade:54,5" *)
    reg s32_val_n9;
    (* src = "src/sreg.spade:54,5" *)
    reg s32_val_n10;
    (* src = "src/sreg.spade:54,5" *)
    reg s32_val_n11;
    (* src = "src/sreg.spade:54,5" *)
    reg s32_val_n12;
    (* src = "src/sreg.spade:54,5" *)
    reg s32_val_n13;
    (* src = "src/sreg.spade:54,5" *)
    reg s32_val_n14;
    (* src = "src/sreg.spade:56,5" *)
    reg \s33_val ;
    (* src = "src/sreg.spade:56,5" *)
    reg s33_val_n1;
    (* src = "src/sreg.spade:56,5" *)
    reg s33_val_n2;
    (* src = "src/sreg.spade:56,5" *)
    reg s33_val_n3;
    (* src = "src/sreg.spade:56,5" *)
    reg s33_val_n4;
    (* src = "src/sreg.spade:56,5" *)
    reg s33_val_n5;
    (* src = "src/sreg.spade:56,5" *)
    reg s33_val_n6;
    (* src = "src/sreg.spade:56,5" *)
    reg s33_val_n7;
    (* src = "src/sreg.spade:56,5" *)
    reg s33_val_n8;
    (* src = "src/sreg.spade:56,5" *)
    reg s33_val_n9;
    (* src = "src/sreg.spade:56,5" *)
    reg s33_val_n10;
    (* src = "src/sreg.spade:56,5" *)
    reg s33_val_n11;
    (* src = "src/sreg.spade:56,5" *)
    reg s33_val_n12;
    (* src = "src/sreg.spade:56,5" *)
    reg s33_val_n13;
    (* src = "src/sreg.spade:56,5" *)
    reg s33_val_n14;
    (* src = "src/sreg.spade:56,5" *)
    reg s33_val_n15;
    (* src = "src/sreg.spade:56,5" *)
    reg \s34_val ;
    (* src = "src/sreg.spade:56,5" *)
    reg s34_val_n1;
    (* src = "src/sreg.spade:56,5" *)
    reg s34_val_n2;
    (* src = "src/sreg.spade:56,5" *)
    reg s34_val_n3;
    (* src = "src/sreg.spade:56,5" *)
    reg s34_val_n4;
    (* src = "src/sreg.spade:56,5" *)
    reg s34_val_n5;
    (* src = "src/sreg.spade:56,5" *)
    reg s34_val_n6;
    (* src = "src/sreg.spade:56,5" *)
    reg s34_val_n7;
    (* src = "src/sreg.spade:56,5" *)
    reg s34_val_n8;
    (* src = "src/sreg.spade:56,5" *)
    reg s34_val_n9;
    (* src = "src/sreg.spade:56,5" *)
    reg s34_val_n10;
    (* src = "src/sreg.spade:56,5" *)
    reg s34_val_n11;
    (* src = "src/sreg.spade:56,5" *)
    reg s34_val_n12;
    (* src = "src/sreg.spade:56,5" *)
    reg s34_val_n13;
    (* src = "src/sreg.spade:56,5" *)
    reg s34_val_n14;
    (* src = "src/sreg.spade:56,5" *)
    reg s34_val_n15;
    (* src = "src/sreg.spade:58,5" *)
    reg \s35_val ;
    (* src = "src/sreg.spade:58,5" *)
    reg s35_val_n1;
    (* src = "src/sreg.spade:58,5" *)
    reg s35_val_n2;
    (* src = "src/sreg.spade:58,5" *)
    reg s35_val_n3;
    (* src = "src/sreg.spade:58,5" *)
    reg s35_val_n4;
    (* src = "src/sreg.spade:58,5" *)
    reg s35_val_n5;
    (* src = "src/sreg.spade:58,5" *)
    reg s35_val_n6;
    (* src = "src/sreg.spade:58,5" *)
    reg s35_val_n7;
    (* src = "src/sreg.spade:58,5" *)
    reg s35_val_n8;
    (* src = "src/sreg.spade:58,5" *)
    reg s35_val_n9;
    (* src = "src/sreg.spade:58,5" *)
    reg s35_val_n10;
    (* src = "src/sreg.spade:58,5" *)
    reg s35_val_n11;
    (* src = "src/sreg.spade:58,5" *)
    reg s35_val_n12;
    (* src = "src/sreg.spade:58,5" *)
    reg s35_val_n13;
    (* src = "src/sreg.spade:58,5" *)
    reg s35_val_n14;
    (* src = "src/sreg.spade:58,5" *)
    reg s35_val_n15;
    (* src = "src/sreg.spade:58,5" *)
    reg s35_val_n16;
    (* src = "src/sreg.spade:58,5" *)
    reg \s36_val ;
    (* src = "src/sreg.spade:58,5" *)
    reg s36_val_n1;
    (* src = "src/sreg.spade:58,5" *)
    reg s36_val_n2;
    (* src = "src/sreg.spade:58,5" *)
    reg s36_val_n3;
    (* src = "src/sreg.spade:58,5" *)
    reg s36_val_n4;
    (* src = "src/sreg.spade:58,5" *)
    reg s36_val_n5;
    (* src = "src/sreg.spade:58,5" *)
    reg s36_val_n6;
    (* src = "src/sreg.spade:58,5" *)
    reg s36_val_n7;
    (* src = "src/sreg.spade:58,5" *)
    reg s36_val_n8;
    (* src = "src/sreg.spade:58,5" *)
    reg s36_val_n9;
    (* src = "src/sreg.spade:58,5" *)
    reg s36_val_n10;
    (* src = "src/sreg.spade:58,5" *)
    reg s36_val_n11;
    (* src = "src/sreg.spade:58,5" *)
    reg s36_val_n12;
    (* src = "src/sreg.spade:58,5" *)
    reg s36_val_n13;
    (* src = "src/sreg.spade:58,5" *)
    reg s36_val_n14;
    (* src = "src/sreg.spade:58,5" *)
    reg s36_val_n15;
    (* src = "src/sreg.spade:58,5" *)
    reg s36_val_n16;
    (* src = "src/sreg.spade:60,5" *)
    reg \s37_val ;
    (* src = "src/sreg.spade:60,5" *)
    reg s37_val_n1;
    (* src = "src/sreg.spade:60,5" *)
    reg s37_val_n2;
    (* src = "src/sreg.spade:60,5" *)
    reg s37_val_n3;
    (* src = "src/sreg.spade:60,5" *)
    reg s37_val_n4;
    (* src = "src/sreg.spade:60,5" *)
    reg s37_val_n5;
    (* src = "src/sreg.spade:60,5" *)
    reg s37_val_n6;
    (* src = "src/sreg.spade:60,5" *)
    reg s37_val_n7;
    (* src = "src/sreg.spade:60,5" *)
    reg s37_val_n8;
    (* src = "src/sreg.spade:60,5" *)
    reg s37_val_n9;
    (* src = "src/sreg.spade:60,5" *)
    reg s37_val_n10;
    (* src = "src/sreg.spade:60,5" *)
    reg s37_val_n11;
    (* src = "src/sreg.spade:60,5" *)
    reg s37_val_n12;
    (* src = "src/sreg.spade:60,5" *)
    reg s37_val_n13;
    (* src = "src/sreg.spade:60,5" *)
    reg s37_val_n14;
    (* src = "src/sreg.spade:60,5" *)
    reg s37_val_n15;
    (* src = "src/sreg.spade:60,5" *)
    reg s37_val_n16;
    (* src = "src/sreg.spade:60,5" *)
    reg s37_val_n17;
    (* src = "src/sreg.spade:60,5" *)
    reg \s38_val ;
    (* src = "src/sreg.spade:60,5" *)
    reg s38_val_n1;
    (* src = "src/sreg.spade:60,5" *)
    reg s38_val_n2;
    (* src = "src/sreg.spade:60,5" *)
    reg s38_val_n3;
    (* src = "src/sreg.spade:60,5" *)
    reg s38_val_n4;
    (* src = "src/sreg.spade:60,5" *)
    reg s38_val_n5;
    (* src = "src/sreg.spade:60,5" *)
    reg s38_val_n6;
    (* src = "src/sreg.spade:60,5" *)
    reg s38_val_n7;
    (* src = "src/sreg.spade:60,5" *)
    reg s38_val_n8;
    (* src = "src/sreg.spade:60,5" *)
    reg s38_val_n9;
    (* src = "src/sreg.spade:60,5" *)
    reg s38_val_n10;
    (* src = "src/sreg.spade:60,5" *)
    reg s38_val_n11;
    (* src = "src/sreg.spade:60,5" *)
    reg s38_val_n12;
    (* src = "src/sreg.spade:60,5" *)
    reg s38_val_n13;
    (* src = "src/sreg.spade:60,5" *)
    reg s38_val_n14;
    (* src = "src/sreg.spade:60,5" *)
    reg s38_val_n15;
    (* src = "src/sreg.spade:60,5" *)
    reg s38_val_n16;
    (* src = "src/sreg.spade:60,5" *)
    reg s38_val_n17;
    (* src = "src/sreg.spade:62,5" *)
    reg \s39_val ;
    (* src = "src/sreg.spade:62,5" *)
    reg s39_val_n1;
    (* src = "src/sreg.spade:62,5" *)
    reg s39_val_n2;
    (* src = "src/sreg.spade:62,5" *)
    reg s39_val_n3;
    (* src = "src/sreg.spade:62,5" *)
    reg s39_val_n4;
    (* src = "src/sreg.spade:62,5" *)
    reg s39_val_n5;
    (* src = "src/sreg.spade:62,5" *)
    reg s39_val_n6;
    (* src = "src/sreg.spade:62,5" *)
    reg s39_val_n7;
    (* src = "src/sreg.spade:62,5" *)
    reg s39_val_n8;
    (* src = "src/sreg.spade:62,5" *)
    reg s39_val_n9;
    (* src = "src/sreg.spade:62,5" *)
    reg s39_val_n10;
    (* src = "src/sreg.spade:62,5" *)
    reg s39_val_n11;
    (* src = "src/sreg.spade:62,5" *)
    reg s39_val_n12;
    (* src = "src/sreg.spade:62,5" *)
    reg s39_val_n13;
    (* src = "src/sreg.spade:62,5" *)
    reg s39_val_n14;
    (* src = "src/sreg.spade:62,5" *)
    reg s39_val_n15;
    (* src = "src/sreg.spade:62,5" *)
    reg s39_val_n16;
    (* src = "src/sreg.spade:62,5" *)
    reg s39_val_n17;
    (* src = "src/sreg.spade:62,5" *)
    reg s39_val_n18;
    (* src = "src/sreg.spade:62,5" *)
    reg \s40_val ;
    (* src = "src/sreg.spade:62,5" *)
    reg s40_val_n1;
    (* src = "src/sreg.spade:62,5" *)
    reg s40_val_n2;
    (* src = "src/sreg.spade:62,5" *)
    reg s40_val_n3;
    (* src = "src/sreg.spade:62,5" *)
    reg s40_val_n4;
    (* src = "src/sreg.spade:62,5" *)
    reg s40_val_n5;
    (* src = "src/sreg.spade:62,5" *)
    reg s40_val_n6;
    (* src = "src/sreg.spade:62,5" *)
    reg s40_val_n7;
    (* src = "src/sreg.spade:62,5" *)
    reg s40_val_n8;
    (* src = "src/sreg.spade:62,5" *)
    reg s40_val_n9;
    (* src = "src/sreg.spade:62,5" *)
    reg s40_val_n10;
    (* src = "src/sreg.spade:62,5" *)
    reg s40_val_n11;
    (* src = "src/sreg.spade:62,5" *)
    reg s40_val_n12;
    (* src = "src/sreg.spade:62,5" *)
    reg s40_val_n13;
    (* src = "src/sreg.spade:62,5" *)
    reg s40_val_n14;
    (* src = "src/sreg.spade:62,5" *)
    reg s40_val_n15;
    (* src = "src/sreg.spade:62,5" *)
    reg s40_val_n16;
    (* src = "src/sreg.spade:62,5" *)
    reg s40_val_n17;
    (* src = "src/sreg.spade:62,5" *)
    reg s40_val_n18;
    (* src = "src/sreg.spade:64,5" *)
    reg \s41_val ;
    (* src = "src/sreg.spade:64,5" *)
    reg s41_val_n1;
    (* src = "src/sreg.spade:64,5" *)
    reg s41_val_n2;
    (* src = "src/sreg.spade:64,5" *)
    reg s41_val_n3;
    (* src = "src/sreg.spade:64,5" *)
    reg s41_val_n4;
    (* src = "src/sreg.spade:64,5" *)
    reg s41_val_n5;
    (* src = "src/sreg.spade:64,5" *)
    reg s41_val_n6;
    (* src = "src/sreg.spade:64,5" *)
    reg s41_val_n7;
    (* src = "src/sreg.spade:64,5" *)
    reg s41_val_n8;
    (* src = "src/sreg.spade:64,5" *)
    reg s41_val_n9;
    (* src = "src/sreg.spade:64,5" *)
    reg s41_val_n10;
    (* src = "src/sreg.spade:64,5" *)
    reg s41_val_n11;
    (* src = "src/sreg.spade:64,5" *)
    reg s41_val_n12;
    (* src = "src/sreg.spade:64,5" *)
    reg s41_val_n13;
    (* src = "src/sreg.spade:64,5" *)
    reg s41_val_n14;
    (* src = "src/sreg.spade:64,5" *)
    reg s41_val_n15;
    (* src = "src/sreg.spade:64,5" *)
    reg s41_val_n16;
    (* src = "src/sreg.spade:64,5" *)
    reg s41_val_n17;
    (* src = "src/sreg.spade:64,5" *)
    reg s41_val_n18;
    (* src = "src/sreg.spade:64,5" *)
    reg s41_val_n19;
    (* src = "src/sreg.spade:64,5" *)
    reg \s42_val ;
    (* src = "src/sreg.spade:64,5" *)
    reg s42_val_n1;
    (* src = "src/sreg.spade:64,5" *)
    reg s42_val_n2;
    (* src = "src/sreg.spade:64,5" *)
    reg s42_val_n3;
    (* src = "src/sreg.spade:64,5" *)
    reg s42_val_n4;
    (* src = "src/sreg.spade:64,5" *)
    reg s42_val_n5;
    (* src = "src/sreg.spade:64,5" *)
    reg s42_val_n6;
    (* src = "src/sreg.spade:64,5" *)
    reg s42_val_n7;
    (* src = "src/sreg.spade:64,5" *)
    reg s42_val_n8;
    (* src = "src/sreg.spade:64,5" *)
    reg s42_val_n9;
    (* src = "src/sreg.spade:64,5" *)
    reg s42_val_n10;
    (* src = "src/sreg.spade:64,5" *)
    reg s42_val_n11;
    (* src = "src/sreg.spade:64,5" *)
    reg s42_val_n12;
    (* src = "src/sreg.spade:64,5" *)
    reg s42_val_n13;
    (* src = "src/sreg.spade:64,5" *)
    reg s42_val_n14;
    (* src = "src/sreg.spade:64,5" *)
    reg s42_val_n15;
    (* src = "src/sreg.spade:64,5" *)
    reg s42_val_n16;
    (* src = "src/sreg.spade:64,5" *)
    reg s42_val_n17;
    (* src = "src/sreg.spade:64,5" *)
    reg s42_val_n18;
    (* src = "src/sreg.spade:64,5" *)
    reg s42_val_n19;
    (* src = "src/sreg.spade:66,5" *)
    reg \s43_val ;
    (* src = "src/sreg.spade:66,5" *)
    reg s43_val_n1;
    (* src = "src/sreg.spade:66,5" *)
    reg s43_val_n2;
    (* src = "src/sreg.spade:66,5" *)
    reg s43_val_n3;
    (* src = "src/sreg.spade:66,5" *)
    reg s43_val_n4;
    (* src = "src/sreg.spade:66,5" *)
    reg s43_val_n5;
    (* src = "src/sreg.spade:66,5" *)
    reg s43_val_n6;
    (* src = "src/sreg.spade:66,5" *)
    reg s43_val_n7;
    (* src = "src/sreg.spade:66,5" *)
    reg s43_val_n8;
    (* src = "src/sreg.spade:66,5" *)
    reg s43_val_n9;
    (* src = "src/sreg.spade:66,5" *)
    reg s43_val_n10;
    (* src = "src/sreg.spade:66,5" *)
    reg s43_val_n11;
    (* src = "src/sreg.spade:66,5" *)
    reg s43_val_n12;
    (* src = "src/sreg.spade:66,5" *)
    reg s43_val_n13;
    (* src = "src/sreg.spade:66,5" *)
    reg s43_val_n14;
    (* src = "src/sreg.spade:66,5" *)
    reg s43_val_n15;
    (* src = "src/sreg.spade:66,5" *)
    reg s43_val_n16;
    (* src = "src/sreg.spade:66,5" *)
    reg s43_val_n17;
    (* src = "src/sreg.spade:66,5" *)
    reg s43_val_n18;
    (* src = "src/sreg.spade:66,5" *)
    reg s43_val_n19;
    (* src = "src/sreg.spade:66,5" *)
    reg s43_val_n20;
    (* src = "src/sreg.spade:66,5" *)
    reg \s44_val ;
    (* src = "src/sreg.spade:66,5" *)
    reg s44_val_n1;
    (* src = "src/sreg.spade:66,5" *)
    reg s44_val_n2;
    (* src = "src/sreg.spade:66,5" *)
    reg s44_val_n3;
    (* src = "src/sreg.spade:66,5" *)
    reg s44_val_n4;
    (* src = "src/sreg.spade:66,5" *)
    reg s44_val_n5;
    (* src = "src/sreg.spade:66,5" *)
    reg s44_val_n6;
    (* src = "src/sreg.spade:66,5" *)
    reg s44_val_n7;
    (* src = "src/sreg.spade:66,5" *)
    reg s44_val_n8;
    (* src = "src/sreg.spade:66,5" *)
    reg s44_val_n9;
    (* src = "src/sreg.spade:66,5" *)
    reg s44_val_n10;
    (* src = "src/sreg.spade:66,5" *)
    reg s44_val_n11;
    (* src = "src/sreg.spade:66,5" *)
    reg s44_val_n12;
    (* src = "src/sreg.spade:66,5" *)
    reg s44_val_n13;
    (* src = "src/sreg.spade:66,5" *)
    reg s44_val_n14;
    (* src = "src/sreg.spade:66,5" *)
    reg s44_val_n15;
    (* src = "src/sreg.spade:66,5" *)
    reg s44_val_n16;
    (* src = "src/sreg.spade:66,5" *)
    reg s44_val_n17;
    (* src = "src/sreg.spade:66,5" *)
    reg s44_val_n18;
    (* src = "src/sreg.spade:66,5" *)
    reg s44_val_n19;
    (* src = "src/sreg.spade:66,5" *)
    reg s44_val_n20;
    (* src = "src/sreg.spade:68,5" *)
    reg \s45_val ;
    (* src = "src/sreg.spade:68,5" *)
    reg s45_val_n1;
    (* src = "src/sreg.spade:68,5" *)
    reg s45_val_n2;
    (* src = "src/sreg.spade:68,5" *)
    reg s45_val_n3;
    (* src = "src/sreg.spade:68,5" *)
    reg s45_val_n4;
    (* src = "src/sreg.spade:68,5" *)
    reg s45_val_n5;
    (* src = "src/sreg.spade:68,5" *)
    reg s45_val_n6;
    (* src = "src/sreg.spade:68,5" *)
    reg s45_val_n7;
    (* src = "src/sreg.spade:68,5" *)
    reg s45_val_n8;
    (* src = "src/sreg.spade:68,5" *)
    reg s45_val_n9;
    (* src = "src/sreg.spade:68,5" *)
    reg s45_val_n10;
    (* src = "src/sreg.spade:68,5" *)
    reg s45_val_n11;
    (* src = "src/sreg.spade:68,5" *)
    reg s45_val_n12;
    (* src = "src/sreg.spade:68,5" *)
    reg s45_val_n13;
    (* src = "src/sreg.spade:68,5" *)
    reg s45_val_n14;
    (* src = "src/sreg.spade:68,5" *)
    reg s45_val_n15;
    (* src = "src/sreg.spade:68,5" *)
    reg s45_val_n16;
    (* src = "src/sreg.spade:68,5" *)
    reg s45_val_n17;
    (* src = "src/sreg.spade:68,5" *)
    reg s45_val_n18;
    (* src = "src/sreg.spade:68,5" *)
    reg s45_val_n19;
    (* src = "src/sreg.spade:68,5" *)
    reg s45_val_n20;
    (* src = "src/sreg.spade:68,5" *)
    reg s45_val_n21;
    (* src = "src/sreg.spade:68,5" *)
    reg \s46_val ;
    (* src = "src/sreg.spade:68,5" *)
    reg s46_val_n1;
    (* src = "src/sreg.spade:68,5" *)
    reg s46_val_n2;
    (* src = "src/sreg.spade:68,5" *)
    reg s46_val_n3;
    (* src = "src/sreg.spade:68,5" *)
    reg s46_val_n4;
    (* src = "src/sreg.spade:68,5" *)
    reg s46_val_n5;
    (* src = "src/sreg.spade:68,5" *)
    reg s46_val_n6;
    (* src = "src/sreg.spade:68,5" *)
    reg s46_val_n7;
    (* src = "src/sreg.spade:68,5" *)
    reg s46_val_n8;
    (* src = "src/sreg.spade:68,5" *)
    reg s46_val_n9;
    (* src = "src/sreg.spade:68,5" *)
    reg s46_val_n10;
    (* src = "src/sreg.spade:68,5" *)
    reg s46_val_n11;
    (* src = "src/sreg.spade:68,5" *)
    reg s46_val_n12;
    (* src = "src/sreg.spade:68,5" *)
    reg s46_val_n13;
    (* src = "src/sreg.spade:68,5" *)
    reg s46_val_n14;
    (* src = "src/sreg.spade:68,5" *)
    reg s46_val_n15;
    (* src = "src/sreg.spade:68,5" *)
    reg s46_val_n16;
    (* src = "src/sreg.spade:68,5" *)
    reg s46_val_n17;
    (* src = "src/sreg.spade:68,5" *)
    reg s46_val_n18;
    (* src = "src/sreg.spade:68,5" *)
    reg s46_val_n19;
    (* src = "src/sreg.spade:68,5" *)
    reg s46_val_n20;
    (* src = "src/sreg.spade:68,5" *)
    reg s46_val_n21;
    (* src = "src/sreg.spade:70,5" *)
    reg \s47_val ;
    (* src = "src/sreg.spade:70,5" *)
    reg s47_val_n1;
    (* src = "src/sreg.spade:70,5" *)
    reg s47_val_n2;
    (* src = "src/sreg.spade:70,5" *)
    reg s47_val_n3;
    (* src = "src/sreg.spade:70,5" *)
    reg s47_val_n4;
    (* src = "src/sreg.spade:70,5" *)
    reg s47_val_n5;
    (* src = "src/sreg.spade:70,5" *)
    reg s47_val_n6;
    (* src = "src/sreg.spade:70,5" *)
    reg s47_val_n7;
    (* src = "src/sreg.spade:70,5" *)
    reg s47_val_n8;
    (* src = "src/sreg.spade:70,5" *)
    reg s47_val_n9;
    (* src = "src/sreg.spade:70,5" *)
    reg s47_val_n10;
    (* src = "src/sreg.spade:70,5" *)
    reg s47_val_n11;
    (* src = "src/sreg.spade:70,5" *)
    reg s47_val_n12;
    (* src = "src/sreg.spade:70,5" *)
    reg s47_val_n13;
    (* src = "src/sreg.spade:70,5" *)
    reg s47_val_n14;
    (* src = "src/sreg.spade:70,5" *)
    reg s47_val_n15;
    (* src = "src/sreg.spade:70,5" *)
    reg s47_val_n16;
    (* src = "src/sreg.spade:70,5" *)
    reg s47_val_n17;
    (* src = "src/sreg.spade:70,5" *)
    reg s47_val_n18;
    (* src = "src/sreg.spade:70,5" *)
    reg s47_val_n19;
    (* src = "src/sreg.spade:70,5" *)
    reg s47_val_n20;
    (* src = "src/sreg.spade:70,5" *)
    reg s47_val_n21;
    (* src = "src/sreg.spade:70,5" *)
    reg s47_val_n22;
    (* src = "src/sreg.spade:70,5" *)
    reg \s48_val ;
    (* src = "src/sreg.spade:70,5" *)
    reg s48_val_n1;
    (* src = "src/sreg.spade:70,5" *)
    reg s48_val_n2;
    (* src = "src/sreg.spade:70,5" *)
    reg s48_val_n3;
    (* src = "src/sreg.spade:70,5" *)
    reg s48_val_n4;
    (* src = "src/sreg.spade:70,5" *)
    reg s48_val_n5;
    (* src = "src/sreg.spade:70,5" *)
    reg s48_val_n6;
    (* src = "src/sreg.spade:70,5" *)
    reg s48_val_n7;
    (* src = "src/sreg.spade:70,5" *)
    reg s48_val_n8;
    (* src = "src/sreg.spade:70,5" *)
    reg s48_val_n9;
    (* src = "src/sreg.spade:70,5" *)
    reg s48_val_n10;
    (* src = "src/sreg.spade:70,5" *)
    reg s48_val_n11;
    (* src = "src/sreg.spade:70,5" *)
    reg s48_val_n12;
    (* src = "src/sreg.spade:70,5" *)
    reg s48_val_n13;
    (* src = "src/sreg.spade:70,5" *)
    reg s48_val_n14;
    (* src = "src/sreg.spade:70,5" *)
    reg s48_val_n15;
    (* src = "src/sreg.spade:70,5" *)
    reg s48_val_n16;
    (* src = "src/sreg.spade:70,5" *)
    reg s48_val_n17;
    (* src = "src/sreg.spade:70,5" *)
    reg s48_val_n18;
    (* src = "src/sreg.spade:70,5" *)
    reg s48_val_n19;
    (* src = "src/sreg.spade:70,5" *)
    reg s48_val_n20;
    (* src = "src/sreg.spade:70,5" *)
    reg s48_val_n21;
    (* src = "src/sreg.spade:70,5" *)
    reg s48_val_n22;
    (* src = "src/sreg.spade:72,5" *)
    reg \s49_val ;
    (* src = "src/sreg.spade:72,5" *)
    reg s49_val_n1;
    (* src = "src/sreg.spade:72,5" *)
    reg s49_val_n2;
    (* src = "src/sreg.spade:72,5" *)
    reg s49_val_n3;
    (* src = "src/sreg.spade:72,5" *)
    reg s49_val_n4;
    (* src = "src/sreg.spade:72,5" *)
    reg s49_val_n5;
    (* src = "src/sreg.spade:72,5" *)
    reg s49_val_n6;
    (* src = "src/sreg.spade:72,5" *)
    reg s49_val_n7;
    (* src = "src/sreg.spade:72,5" *)
    reg s49_val_n8;
    (* src = "src/sreg.spade:72,5" *)
    reg s49_val_n9;
    (* src = "src/sreg.spade:72,5" *)
    reg s49_val_n10;
    (* src = "src/sreg.spade:72,5" *)
    reg s49_val_n11;
    (* src = "src/sreg.spade:72,5" *)
    reg s49_val_n12;
    (* src = "src/sreg.spade:72,5" *)
    reg s49_val_n13;
    (* src = "src/sreg.spade:72,5" *)
    reg s49_val_n14;
    (* src = "src/sreg.spade:72,5" *)
    reg s49_val_n15;
    (* src = "src/sreg.spade:72,5" *)
    reg s49_val_n16;
    (* src = "src/sreg.spade:72,5" *)
    reg s49_val_n17;
    (* src = "src/sreg.spade:72,5" *)
    reg s49_val_n18;
    (* src = "src/sreg.spade:72,5" *)
    reg s49_val_n19;
    (* src = "src/sreg.spade:72,5" *)
    reg s49_val_n20;
    (* src = "src/sreg.spade:72,5" *)
    reg s49_val_n21;
    (* src = "src/sreg.spade:72,5" *)
    reg s49_val_n22;
    (* src = "src/sreg.spade:72,5" *)
    reg s49_val_n23;
    (* src = "src/sreg.spade:72,5" *)
    reg \s50_val ;
    (* src = "src/sreg.spade:72,5" *)
    reg s50_val_n1;
    (* src = "src/sreg.spade:72,5" *)
    reg s50_val_n2;
    (* src = "src/sreg.spade:72,5" *)
    reg s50_val_n3;
    (* src = "src/sreg.spade:72,5" *)
    reg s50_val_n4;
    (* src = "src/sreg.spade:72,5" *)
    reg s50_val_n5;
    (* src = "src/sreg.spade:72,5" *)
    reg s50_val_n6;
    (* src = "src/sreg.spade:72,5" *)
    reg s50_val_n7;
    (* src = "src/sreg.spade:72,5" *)
    reg s50_val_n8;
    (* src = "src/sreg.spade:72,5" *)
    reg s50_val_n9;
    (* src = "src/sreg.spade:72,5" *)
    reg s50_val_n10;
    (* src = "src/sreg.spade:72,5" *)
    reg s50_val_n11;
    (* src = "src/sreg.spade:72,5" *)
    reg s50_val_n12;
    (* src = "src/sreg.spade:72,5" *)
    reg s50_val_n13;
    (* src = "src/sreg.spade:72,5" *)
    reg s50_val_n14;
    (* src = "src/sreg.spade:72,5" *)
    reg s50_val_n15;
    (* src = "src/sreg.spade:72,5" *)
    reg s50_val_n16;
    (* src = "src/sreg.spade:72,5" *)
    reg s50_val_n17;
    (* src = "src/sreg.spade:72,5" *)
    reg s50_val_n18;
    (* src = "src/sreg.spade:72,5" *)
    reg s50_val_n19;
    (* src = "src/sreg.spade:72,5" *)
    reg s50_val_n20;
    (* src = "src/sreg.spade:72,5" *)
    reg s50_val_n21;
    (* src = "src/sreg.spade:72,5" *)
    reg s50_val_n22;
    (* src = "src/sreg.spade:72,5" *)
    reg s50_val_n23;
    (* src = "src/sreg.spade:74,5" *)
    reg \s51_val ;
    (* src = "src/sreg.spade:74,5" *)
    reg s51_val_n1;
    (* src = "src/sreg.spade:74,5" *)
    reg s51_val_n2;
    (* src = "src/sreg.spade:74,5" *)
    reg s51_val_n3;
    (* src = "src/sreg.spade:74,5" *)
    reg s51_val_n4;
    (* src = "src/sreg.spade:74,5" *)
    reg s51_val_n5;
    (* src = "src/sreg.spade:74,5" *)
    reg s51_val_n6;
    (* src = "src/sreg.spade:74,5" *)
    reg s51_val_n7;
    (* src = "src/sreg.spade:74,5" *)
    reg s51_val_n8;
    (* src = "src/sreg.spade:74,5" *)
    reg s51_val_n9;
    (* src = "src/sreg.spade:74,5" *)
    reg s51_val_n10;
    (* src = "src/sreg.spade:74,5" *)
    reg s51_val_n11;
    (* src = "src/sreg.spade:74,5" *)
    reg s51_val_n12;
    (* src = "src/sreg.spade:74,5" *)
    reg s51_val_n13;
    (* src = "src/sreg.spade:74,5" *)
    reg s51_val_n14;
    (* src = "src/sreg.spade:74,5" *)
    reg s51_val_n15;
    (* src = "src/sreg.spade:74,5" *)
    reg s51_val_n16;
    (* src = "src/sreg.spade:74,5" *)
    reg s51_val_n17;
    (* src = "src/sreg.spade:74,5" *)
    reg s51_val_n18;
    (* src = "src/sreg.spade:74,5" *)
    reg s51_val_n19;
    (* src = "src/sreg.spade:74,5" *)
    reg s51_val_n20;
    (* src = "src/sreg.spade:74,5" *)
    reg s51_val_n21;
    (* src = "src/sreg.spade:74,5" *)
    reg s51_val_n22;
    (* src = "src/sreg.spade:74,5" *)
    reg s51_val_n23;
    (* src = "src/sreg.spade:74,5" *)
    reg s51_val_n24;
    (* src = "src/sreg.spade:74,5" *)
    reg \s52_val ;
    (* src = "src/sreg.spade:74,5" *)
    reg s52_val_n1;
    (* src = "src/sreg.spade:74,5" *)
    reg s52_val_n2;
    (* src = "src/sreg.spade:74,5" *)
    reg s52_val_n3;
    (* src = "src/sreg.spade:74,5" *)
    reg s52_val_n4;
    (* src = "src/sreg.spade:74,5" *)
    reg s52_val_n5;
    (* src = "src/sreg.spade:74,5" *)
    reg s52_val_n6;
    (* src = "src/sreg.spade:74,5" *)
    reg s52_val_n7;
    (* src = "src/sreg.spade:74,5" *)
    reg s52_val_n8;
    (* src = "src/sreg.spade:74,5" *)
    reg s52_val_n9;
    (* src = "src/sreg.spade:74,5" *)
    reg s52_val_n10;
    (* src = "src/sreg.spade:74,5" *)
    reg s52_val_n11;
    (* src = "src/sreg.spade:74,5" *)
    reg s52_val_n12;
    (* src = "src/sreg.spade:74,5" *)
    reg s52_val_n13;
    (* src = "src/sreg.spade:74,5" *)
    reg s52_val_n14;
    (* src = "src/sreg.spade:74,5" *)
    reg s52_val_n15;
    (* src = "src/sreg.spade:74,5" *)
    reg s52_val_n16;
    (* src = "src/sreg.spade:74,5" *)
    reg s52_val_n17;
    (* src = "src/sreg.spade:74,5" *)
    reg s52_val_n18;
    (* src = "src/sreg.spade:74,5" *)
    reg s52_val_n19;
    (* src = "src/sreg.spade:74,5" *)
    reg s52_val_n20;
    (* src = "src/sreg.spade:74,5" *)
    reg s52_val_n21;
    (* src = "src/sreg.spade:74,5" *)
    reg s52_val_n22;
    (* src = "src/sreg.spade:74,5" *)
    reg s52_val_n23;
    (* src = "src/sreg.spade:74,5" *)
    reg s52_val_n24;
    (* src = "src/sreg.spade:76,5" *)
    reg \s53_val ;
    (* src = "src/sreg.spade:76,5" *)
    reg s53_val_n1;
    (* src = "src/sreg.spade:76,5" *)
    reg s53_val_n2;
    (* src = "src/sreg.spade:76,5" *)
    reg s53_val_n3;
    (* src = "src/sreg.spade:76,5" *)
    reg s53_val_n4;
    (* src = "src/sreg.spade:76,5" *)
    reg s53_val_n5;
    (* src = "src/sreg.spade:76,5" *)
    reg s53_val_n6;
    (* src = "src/sreg.spade:76,5" *)
    reg s53_val_n7;
    (* src = "src/sreg.spade:76,5" *)
    reg s53_val_n8;
    (* src = "src/sreg.spade:76,5" *)
    reg s53_val_n9;
    (* src = "src/sreg.spade:76,5" *)
    reg s53_val_n10;
    (* src = "src/sreg.spade:76,5" *)
    reg s53_val_n11;
    (* src = "src/sreg.spade:76,5" *)
    reg s53_val_n12;
    (* src = "src/sreg.spade:76,5" *)
    reg s53_val_n13;
    (* src = "src/sreg.spade:76,5" *)
    reg s53_val_n14;
    (* src = "src/sreg.spade:76,5" *)
    reg s53_val_n15;
    (* src = "src/sreg.spade:76,5" *)
    reg s53_val_n16;
    (* src = "src/sreg.spade:76,5" *)
    reg s53_val_n17;
    (* src = "src/sreg.spade:76,5" *)
    reg s53_val_n18;
    (* src = "src/sreg.spade:76,5" *)
    reg s53_val_n19;
    (* src = "src/sreg.spade:76,5" *)
    reg s53_val_n20;
    (* src = "src/sreg.spade:76,5" *)
    reg s53_val_n21;
    (* src = "src/sreg.spade:76,5" *)
    reg s53_val_n22;
    (* src = "src/sreg.spade:76,5" *)
    reg s53_val_n23;
    (* src = "src/sreg.spade:76,5" *)
    reg s53_val_n24;
    (* src = "src/sreg.spade:76,5" *)
    reg s53_val_n25;
    (* src = "src/sreg.spade:76,5" *)
    reg \s54_val ;
    (* src = "src/sreg.spade:76,5" *)
    reg s54_val_n1;
    (* src = "src/sreg.spade:76,5" *)
    reg s54_val_n2;
    (* src = "src/sreg.spade:76,5" *)
    reg s54_val_n3;
    (* src = "src/sreg.spade:76,5" *)
    reg s54_val_n4;
    (* src = "src/sreg.spade:76,5" *)
    reg s54_val_n5;
    (* src = "src/sreg.spade:76,5" *)
    reg s54_val_n6;
    (* src = "src/sreg.spade:76,5" *)
    reg s54_val_n7;
    (* src = "src/sreg.spade:76,5" *)
    reg s54_val_n8;
    (* src = "src/sreg.spade:76,5" *)
    reg s54_val_n9;
    (* src = "src/sreg.spade:76,5" *)
    reg s54_val_n10;
    (* src = "src/sreg.spade:76,5" *)
    reg s54_val_n11;
    (* src = "src/sreg.spade:76,5" *)
    reg s54_val_n12;
    (* src = "src/sreg.spade:76,5" *)
    reg s54_val_n13;
    (* src = "src/sreg.spade:76,5" *)
    reg s54_val_n14;
    (* src = "src/sreg.spade:76,5" *)
    reg s54_val_n15;
    (* src = "src/sreg.spade:76,5" *)
    reg s54_val_n16;
    (* src = "src/sreg.spade:76,5" *)
    reg s54_val_n17;
    (* src = "src/sreg.spade:76,5" *)
    reg s54_val_n18;
    (* src = "src/sreg.spade:76,5" *)
    reg s54_val_n19;
    (* src = "src/sreg.spade:76,5" *)
    reg s54_val_n20;
    (* src = "src/sreg.spade:76,5" *)
    reg s54_val_n21;
    (* src = "src/sreg.spade:76,5" *)
    reg s54_val_n22;
    (* src = "src/sreg.spade:76,5" *)
    reg s54_val_n23;
    (* src = "src/sreg.spade:76,5" *)
    reg s54_val_n24;
    (* src = "src/sreg.spade:76,5" *)
    reg s54_val_n25;
    (* src = "src/sreg.spade:78,5" *)
    reg \s55_val ;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n1;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n2;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n3;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n4;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n5;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n6;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n7;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n8;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n9;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n10;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n11;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n12;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n13;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n14;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n15;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n16;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n17;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n18;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n19;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n20;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n21;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n22;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n23;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n24;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n25;
    (* src = "src/sreg.spade:78,5" *)
    reg s55_val_n26;
    (* src = "src/sreg.spade:78,5" *)
    reg \s56_val ;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n1;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n2;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n3;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n4;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n5;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n6;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n7;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n8;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n9;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n10;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n11;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n12;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n13;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n14;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n15;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n16;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n17;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n18;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n19;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n20;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n21;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n22;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n23;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n24;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n25;
    (* src = "src/sreg.spade:78,5" *)
    reg s56_val_n26;
    (* src = "src/sreg.spade:80,5" *)
    reg \s57_val ;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n1;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n2;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n3;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n4;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n5;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n6;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n7;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n8;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n9;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n10;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n11;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n12;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n13;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n14;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n15;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n16;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n17;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n18;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n19;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n20;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n21;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n22;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n23;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n24;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n25;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n26;
    (* src = "src/sreg.spade:80,5" *)
    reg s57_val_n27;
    (* src = "src/sreg.spade:80,5" *)
    reg \s58_val ;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n1;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n2;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n3;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n4;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n5;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n6;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n7;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n8;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n9;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n10;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n11;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n12;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n13;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n14;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n15;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n16;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n17;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n18;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n19;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n20;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n21;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n22;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n23;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n24;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n25;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n26;
    (* src = "src/sreg.spade:80,5" *)
    reg s58_val_n27;
    (* src = "src/sreg.spade:82,5" *)
    reg \s59_val ;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n1;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n2;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n3;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n4;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n5;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n6;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n7;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n8;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n9;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n10;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n11;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n12;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n13;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n14;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n15;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n16;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n17;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n18;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n19;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n20;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n21;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n22;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n23;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n24;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n25;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n26;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n27;
    (* src = "src/sreg.spade:82,5" *)
    reg s59_val_n28;
    (* src = "src/sreg.spade:82,5" *)
    reg \s60_val ;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n1;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n2;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n3;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n4;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n5;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n6;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n7;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n8;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n9;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n10;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n11;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n12;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n13;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n14;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n15;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n16;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n17;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n18;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n19;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n20;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n21;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n22;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n23;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n24;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n25;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n26;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n27;
    (* src = "src/sreg.spade:82,5" *)
    reg s60_val_n28;
    (* src = "src/sreg.spade:84,5" *)
    reg \s61_val ;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n1;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n2;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n3;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n4;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n5;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n6;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n7;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n8;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n9;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n10;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n11;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n12;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n13;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n14;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n15;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n16;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n17;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n18;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n19;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n20;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n21;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n22;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n23;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n24;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n25;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n26;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n27;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n28;
    (* src = "src/sreg.spade:84,5" *)
    reg s61_val_n29;
    (* src = "src/sreg.spade:84,5" *)
    reg \s62_val ;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n1;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n2;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n3;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n4;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n5;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n6;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n7;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n8;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n9;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n10;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n11;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n12;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n13;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n14;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n15;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n16;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n17;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n18;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n19;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n20;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n21;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n22;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n23;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n24;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n25;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n26;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n27;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n28;
    (* src = "src/sreg.spade:84,5" *)
    reg s62_val_n29;
    (* src = "src/sreg.spade:86,5" *)
    reg \s63_val ;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n1;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n2;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n3;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n4;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n5;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n6;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n7;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n8;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n9;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n10;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n11;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n12;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n13;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n14;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n15;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n16;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n17;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n18;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n19;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n20;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n21;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n22;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n23;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n24;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n25;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n26;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n27;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n28;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n29;
    (* src = "src/sreg.spade:86,5" *)
    reg s63_val_n30;
    (* src = "src/sreg.spade:86,5" *)
    reg \s64_val ;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n1;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n2;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n3;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n4;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n5;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n6;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n7;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n8;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n9;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n10;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n11;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n12;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n13;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n14;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n15;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n16;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n17;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n18;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n19;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n20;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n21;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n22;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n23;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n24;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n25;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n26;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n27;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n28;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n29;
    (* src = "src/sreg.spade:86,5" *)
    reg s64_val_n30;
    (* src = "src/sreg.spade:88,5" *)
    reg \s65_val ;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n1;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n2;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n3;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n4;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n5;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n6;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n7;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n8;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n9;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n10;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n11;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n12;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n13;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n14;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n15;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n16;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n17;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n18;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n19;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n20;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n21;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n22;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n23;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n24;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n25;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n26;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n27;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n28;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n29;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n30;
    (* src = "src/sreg.spade:88,5" *)
    reg s65_val_n31;
    (* src = "src/sreg.spade:88,5" *)
    reg \s66_val ;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n1;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n2;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n3;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n4;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n5;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n6;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n7;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n8;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n9;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n10;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n11;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n12;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n13;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n14;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n15;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n16;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n17;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n18;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n19;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n20;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n21;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n22;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n23;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n24;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n25;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n26;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n27;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n28;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n29;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n30;
    (* src = "src/sreg.spade:88,5" *)
    reg s66_val_n31;
    (* src = "src/sreg.spade:90,5" *)
    reg \s67_val ;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n1;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n2;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n3;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n4;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n5;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n6;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n7;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n8;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n9;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n10;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n11;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n12;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n13;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n14;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n15;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n16;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n17;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n18;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n19;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n20;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n21;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n22;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n23;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n24;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n25;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n26;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n27;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n28;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n29;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n30;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n31;
    (* src = "src/sreg.spade:90,5" *)
    reg s67_val_n32;
    (* src = "src/sreg.spade:90,5" *)
    reg \s68_val ;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n1;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n2;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n3;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n4;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n5;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n6;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n7;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n8;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n9;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n10;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n11;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n12;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n13;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n14;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n15;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n16;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n17;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n18;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n19;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n20;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n21;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n22;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n23;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n24;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n25;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n26;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n27;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n28;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n29;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n30;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n31;
    (* src = "src/sreg.spade:90,5" *)
    reg s68_val_n32;
    (* src = "src/sreg.spade:92,5" *)
    reg \s69_val ;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n1;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n2;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n3;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n4;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n5;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n6;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n7;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n8;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n9;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n10;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n11;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n12;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n13;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n14;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n15;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n16;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n17;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n18;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n19;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n20;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n21;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n22;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n23;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n24;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n25;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n26;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n27;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n28;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n29;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n30;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n31;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n32;
    (* src = "src/sreg.spade:92,5" *)
    reg s69_val_n33;
    (* src = "src/sreg.spade:92,5" *)
    reg \s70_val ;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n1;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n2;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n3;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n4;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n5;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n6;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n7;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n8;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n9;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n10;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n11;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n12;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n13;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n14;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n15;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n16;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n17;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n18;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n19;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n20;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n21;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n22;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n23;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n24;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n25;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n26;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n27;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n28;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n29;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n30;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n31;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n32;
    (* src = "src/sreg.spade:92,5" *)
    reg s70_val_n33;
    (* src = "src/sreg.spade:94,5" *)
    reg \s71_val ;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n1;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n2;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n3;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n4;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n5;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n6;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n7;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n8;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n9;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n10;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n11;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n12;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n13;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n14;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n15;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n16;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n17;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n18;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n19;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n20;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n21;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n22;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n23;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n24;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n25;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n26;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n27;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n28;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n29;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n30;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n31;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n32;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n33;
    (* src = "src/sreg.spade:94,5" *)
    reg s71_val_n34;
    (* src = "src/sreg.spade:94,5" *)
    reg \s72_val ;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n1;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n2;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n3;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n4;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n5;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n6;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n7;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n8;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n9;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n10;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n11;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n12;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n13;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n14;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n15;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n16;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n17;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n18;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n19;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n20;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n21;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n22;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n23;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n24;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n25;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n26;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n27;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n28;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n29;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n30;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n31;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n32;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n33;
    (* src = "src/sreg.spade:94,5" *)
    reg s72_val_n34;
    (* src = "src/sreg.spade:96,5" *)
    reg \s73_val ;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n1;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n2;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n3;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n4;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n5;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n6;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n7;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n8;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n9;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n10;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n11;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n12;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n13;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n14;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n15;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n16;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n17;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n18;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n19;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n20;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n21;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n22;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n23;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n24;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n25;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n26;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n27;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n28;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n29;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n30;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n31;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n32;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n33;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n34;
    (* src = "src/sreg.spade:96,5" *)
    reg s73_val_n35;
    (* src = "src/sreg.spade:96,5" *)
    reg \s74_val ;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n1;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n2;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n3;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n4;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n5;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n6;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n7;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n8;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n9;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n10;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n11;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n12;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n13;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n14;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n15;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n16;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n17;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n18;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n19;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n20;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n21;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n22;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n23;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n24;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n25;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n26;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n27;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n28;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n29;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n30;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n31;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n32;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n33;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n34;
    (* src = "src/sreg.spade:96,5" *)
    reg s74_val_n35;
    (* src = "src/sreg.spade:98,5" *)
    reg \s75_val ;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n1;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n2;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n3;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n4;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n5;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n6;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n7;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n8;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n9;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n10;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n11;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n12;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n13;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n14;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n15;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n16;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n17;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n18;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n19;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n20;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n21;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n22;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n23;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n24;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n25;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n26;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n27;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n28;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n29;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n30;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n31;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n32;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n33;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n34;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n35;
    (* src = "src/sreg.spade:98,5" *)
    reg s75_val_n36;
    (* src = "src/sreg.spade:98,5" *)
    reg \s76_val ;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n1;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n2;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n3;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n4;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n5;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n6;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n7;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n8;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n9;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n10;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n11;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n12;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n13;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n14;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n15;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n16;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n17;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n18;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n19;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n20;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n21;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n22;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n23;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n24;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n25;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n26;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n27;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n28;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n29;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n30;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n31;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n32;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n33;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n34;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n35;
    (* src = "src/sreg.spade:98,5" *)
    reg s76_val_n36;
    (* src = "src/sreg.spade:100,5" *)
    reg \s77_val ;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n1;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n2;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n3;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n4;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n5;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n6;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n7;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n8;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n9;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n10;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n11;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n12;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n13;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n14;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n15;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n16;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n17;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n18;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n19;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n20;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n21;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n22;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n23;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n24;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n25;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n26;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n27;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n28;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n29;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n30;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n31;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n32;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n33;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n34;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n35;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n36;
    (* src = "src/sreg.spade:100,5" *)
    reg s77_val_n37;
    (* src = "src/sreg.spade:100,5" *)
    reg \s78_val ;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n1;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n2;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n3;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n4;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n5;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n6;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n7;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n8;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n9;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n10;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n11;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n12;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n13;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n14;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n15;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n16;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n17;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n18;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n19;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n20;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n21;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n22;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n23;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n24;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n25;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n26;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n27;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n28;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n29;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n30;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n31;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n32;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n33;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n34;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n35;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n36;
    (* src = "src/sreg.spade:100,5" *)
    reg s78_val_n37;
    (* src = "src/sreg.spade:102,5" *)
    reg \s79_val ;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n1;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n2;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n3;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n4;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n5;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n6;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n7;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n8;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n9;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n10;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n11;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n12;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n13;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n14;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n15;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n16;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n17;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n18;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n19;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n20;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n21;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n22;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n23;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n24;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n25;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n26;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n27;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n28;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n29;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n30;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n31;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n32;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n33;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n34;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n35;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n36;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n37;
    (* src = "src/sreg.spade:102,5" *)
    reg s79_val_n38;
    (* src = "src/sreg.spade:102,5" *)
    reg \s80_val ;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n1;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n2;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n3;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n4;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n5;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n6;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n7;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n8;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n9;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n10;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n11;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n12;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n13;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n14;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n15;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n16;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n17;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n18;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n19;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n20;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n21;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n22;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n23;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n24;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n25;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n26;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n27;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n28;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n29;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n30;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n31;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n32;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n33;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n34;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n35;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n36;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n37;
    (* src = "src/sreg.spade:102,5" *)
    reg s80_val_n38;
    (* src = "src/sreg.spade:104,5" *)
    reg \s81_val ;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n1;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n2;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n3;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n4;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n5;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n6;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n7;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n8;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n9;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n10;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n11;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n12;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n13;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n14;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n15;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n16;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n17;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n18;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n19;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n20;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n21;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n22;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n23;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n24;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n25;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n26;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n27;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n28;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n29;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n30;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n31;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n32;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n33;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n34;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n35;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n36;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n37;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n38;
    (* src = "src/sreg.spade:104,5" *)
    reg s81_val_n39;
    (* src = "src/sreg.spade:104,5" *)
    reg \s82_val ;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n1;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n2;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n3;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n4;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n5;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n6;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n7;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n8;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n9;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n10;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n11;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n12;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n13;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n14;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n15;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n16;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n17;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n18;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n19;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n20;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n21;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n22;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n23;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n24;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n25;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n26;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n27;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n28;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n29;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n30;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n31;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n32;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n33;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n34;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n35;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n36;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n37;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n38;
    (* src = "src/sreg.spade:104,5" *)
    reg s82_val_n39;
    (* src = "src/sreg.spade:106,5" *)
    reg \s83_val ;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n1;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n2;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n3;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n4;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n5;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n6;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n7;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n8;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n9;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n10;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n11;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n12;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n13;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n14;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n15;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n16;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n17;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n18;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n19;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n20;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n21;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n22;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n23;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n24;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n25;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n26;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n27;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n28;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n29;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n30;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n31;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n32;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n33;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n34;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n35;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n36;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n37;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n38;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n39;
    (* src = "src/sreg.spade:106,5" *)
    reg s83_val_n40;
    (* src = "src/sreg.spade:106,5" *)
    reg \s84_val ;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n1;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n2;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n3;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n4;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n5;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n6;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n7;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n8;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n9;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n10;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n11;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n12;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n13;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n14;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n15;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n16;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n17;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n18;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n19;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n20;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n21;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n22;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n23;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n24;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n25;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n26;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n27;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n28;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n29;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n30;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n31;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n32;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n33;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n34;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n35;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n36;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n37;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n38;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n39;
    (* src = "src/sreg.spade:106,5" *)
    reg s84_val_n40;
    (* src = "src/sreg.spade:108,5" *)
    reg \s85_val ;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n1;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n2;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n3;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n4;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n5;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n6;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n7;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n8;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n9;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n10;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n11;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n12;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n13;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n14;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n15;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n16;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n17;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n18;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n19;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n20;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n21;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n22;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n23;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n24;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n25;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n26;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n27;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n28;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n29;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n30;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n31;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n32;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n33;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n34;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n35;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n36;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n37;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n38;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n39;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n40;
    (* src = "src/sreg.spade:108,5" *)
    reg s85_val_n41;
    (* src = "src/sreg.spade:108,5" *)
    reg \s86_val ;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n1;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n2;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n3;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n4;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n5;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n6;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n7;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n8;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n9;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n10;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n11;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n12;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n13;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n14;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n15;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n16;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n17;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n18;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n19;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n20;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n21;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n22;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n23;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n24;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n25;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n26;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n27;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n28;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n29;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n30;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n31;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n32;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n33;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n34;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n35;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n36;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n37;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n38;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n39;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n40;
    (* src = "src/sreg.spade:108,5" *)
    reg s86_val_n41;
    (* src = "src/sreg.spade:110,5" *)
    reg \s87_val ;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n1;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n2;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n3;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n4;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n5;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n6;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n7;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n8;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n9;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n10;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n11;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n12;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n13;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n14;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n15;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n16;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n17;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n18;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n19;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n20;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n21;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n22;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n23;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n24;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n25;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n26;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n27;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n28;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n29;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n30;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n31;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n32;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n33;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n34;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n35;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n36;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n37;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n38;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n39;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n40;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n41;
    (* src = "src/sreg.spade:110,5" *)
    reg s87_val_n42;
    (* src = "src/sreg.spade:110,5" *)
    reg \s88_val ;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n1;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n2;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n3;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n4;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n5;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n6;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n7;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n8;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n9;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n10;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n11;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n12;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n13;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n14;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n15;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n16;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n17;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n18;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n19;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n20;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n21;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n22;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n23;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n24;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n25;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n26;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n27;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n28;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n29;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n30;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n31;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n32;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n33;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n34;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n35;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n36;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n37;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n38;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n39;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n40;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n41;
    (* src = "src/sreg.spade:110,5" *)
    reg s88_val_n42;
    (* src = "src/sreg.spade:112,5" *)
    reg \s89_val ;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n1;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n2;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n3;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n4;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n5;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n6;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n7;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n8;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n9;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n10;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n11;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n12;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n13;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n14;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n15;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n16;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n17;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n18;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n19;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n20;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n21;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n22;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n23;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n24;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n25;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n26;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n27;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n28;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n29;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n30;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n31;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n32;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n33;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n34;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n35;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n36;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n37;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n38;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n39;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n40;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n41;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n42;
    (* src = "src/sreg.spade:112,5" *)
    reg s89_val_n43;
    (* src = "src/sreg.spade:112,5" *)
    reg \s90_val ;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n1;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n2;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n3;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n4;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n5;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n6;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n7;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n8;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n9;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n10;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n11;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n12;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n13;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n14;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n15;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n16;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n17;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n18;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n19;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n20;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n21;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n22;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n23;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n24;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n25;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n26;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n27;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n28;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n29;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n30;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n31;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n32;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n33;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n34;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n35;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n36;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n37;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n38;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n39;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n40;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n41;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n42;
    (* src = "src/sreg.spade:112,5" *)
    reg s90_val_n43;
    (* src = "src/sreg.spade:114,5" *)
    reg \s91_val ;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n1;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n2;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n3;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n4;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n5;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n6;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n7;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n8;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n9;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n10;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n11;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n12;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n13;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n14;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n15;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n16;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n17;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n18;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n19;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n20;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n21;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n22;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n23;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n24;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n25;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n26;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n27;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n28;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n29;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n30;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n31;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n32;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n33;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n34;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n35;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n36;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n37;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n38;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n39;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n40;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n41;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n42;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n43;
    (* src = "src/sreg.spade:114,5" *)
    reg s91_val_n44;
    (* src = "src/sreg.spade:114,5" *)
    reg \s92_val ;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n1;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n2;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n3;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n4;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n5;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n6;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n7;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n8;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n9;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n10;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n11;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n12;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n13;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n14;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n15;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n16;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n17;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n18;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n19;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n20;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n21;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n22;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n23;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n24;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n25;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n26;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n27;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n28;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n29;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n30;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n31;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n32;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n33;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n34;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n35;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n36;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n37;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n38;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n39;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n40;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n41;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n42;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n43;
    (* src = "src/sreg.spade:114,5" *)
    reg s92_val_n44;
    (* src = "src/sreg.spade:116,5" *)
    reg \s93_val ;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n1;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n2;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n3;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n4;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n5;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n6;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n7;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n8;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n9;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n10;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n11;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n12;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n13;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n14;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n15;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n16;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n17;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n18;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n19;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n20;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n21;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n22;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n23;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n24;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n25;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n26;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n27;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n28;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n29;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n30;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n31;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n32;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n33;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n34;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n35;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n36;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n37;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n38;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n39;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n40;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n41;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n42;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n43;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n44;
    (* src = "src/sreg.spade:116,5" *)
    reg s93_val_n45;
    (* src = "src/sreg.spade:116,5" *)
    reg \s94_val ;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n1;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n2;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n3;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n4;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n5;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n6;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n7;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n8;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n9;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n10;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n11;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n12;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n13;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n14;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n15;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n16;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n17;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n18;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n19;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n20;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n21;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n22;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n23;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n24;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n25;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n26;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n27;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n28;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n29;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n30;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n31;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n32;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n33;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n34;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n35;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n36;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n37;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n38;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n39;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n40;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n41;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n42;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n43;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n44;
    (* src = "src/sreg.spade:116,5" *)
    reg s94_val_n45;
    (* src = "src/sreg.spade:118,5" *)
    reg \s95_val ;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n1;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n2;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n3;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n4;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n5;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n6;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n7;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n8;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n9;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n10;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n11;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n12;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n13;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n14;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n15;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n16;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n17;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n18;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n19;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n20;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n21;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n22;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n23;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n24;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n25;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n26;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n27;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n28;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n29;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n30;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n31;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n32;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n33;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n34;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n35;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n36;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n37;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n38;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n39;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n40;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n41;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n42;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n43;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n44;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n45;
    (* src = "src/sreg.spade:118,5" *)
    reg s95_val_n46;
    (* src = "src/sreg.spade:118,5" *)
    reg \s96_val ;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n1;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n2;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n3;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n4;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n5;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n6;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n7;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n8;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n9;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n10;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n11;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n12;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n13;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n14;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n15;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n16;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n17;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n18;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n19;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n20;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n21;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n22;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n23;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n24;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n25;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n26;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n27;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n28;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n29;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n30;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n31;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n32;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n33;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n34;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n35;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n36;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n37;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n38;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n39;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n40;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n41;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n42;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n43;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n44;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n45;
    (* src = "src/sreg.spade:118,5" *)
    reg s96_val_n46;
    (* src = "src/sreg.spade:120,5" *)
    reg \s97_val ;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n1;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n2;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n3;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n4;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n5;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n6;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n7;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n8;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n9;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n10;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n11;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n12;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n13;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n14;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n15;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n16;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n17;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n18;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n19;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n20;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n21;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n22;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n23;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n24;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n25;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n26;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n27;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n28;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n29;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n30;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n31;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n32;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n33;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n34;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n35;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n36;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n37;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n38;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n39;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n40;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n41;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n42;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n43;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n44;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n45;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n46;
    (* src = "src/sreg.spade:120,5" *)
    reg s97_val_n47;
    (* src = "src/sreg.spade:120,5" *)
    reg \s98_val ;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n1;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n2;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n3;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n4;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n5;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n6;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n7;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n8;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n9;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n10;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n11;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n12;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n13;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n14;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n15;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n16;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n17;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n18;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n19;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n20;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n21;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n22;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n23;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n24;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n25;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n26;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n27;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n28;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n29;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n30;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n31;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n32;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n33;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n34;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n35;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n36;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n37;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n38;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n39;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n40;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n41;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n42;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n43;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n44;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n45;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n46;
    (* src = "src/sreg.spade:120,5" *)
    reg s98_val_n47;
    (* src = "src/sreg.spade:122,5" *)
    reg \s99_val ;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n1;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n2;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n3;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n4;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n5;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n6;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n7;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n8;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n9;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n10;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n11;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n12;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n13;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n14;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n15;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n16;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n17;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n18;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n19;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n20;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n21;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n22;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n23;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n24;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n25;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n26;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n27;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n28;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n29;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n30;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n31;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n32;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n33;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n34;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n35;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n36;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n37;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n38;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n39;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n40;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n41;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n42;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n43;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n44;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n45;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n46;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n47;
    (* src = "src/sreg.spade:122,5" *)
    reg s99_val_n48;
    (* src = "src/sreg.spade:122,5" *)
    reg \s100_val ;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n1;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n2;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n3;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n4;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n5;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n6;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n7;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n8;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n9;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n10;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n11;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n12;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n13;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n14;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n15;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n16;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n17;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n18;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n19;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n20;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n21;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n22;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n23;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n24;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n25;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n26;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n27;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n28;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n29;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n30;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n31;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n32;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n33;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n34;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n35;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n36;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n37;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n38;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n39;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n40;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n41;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n42;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n43;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n44;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n45;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n46;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n47;
    (* src = "src/sreg.spade:122,5" *)
    reg s100_val_n48;
    (* src = "src/sreg.spade:25,19" *)
    logic val_n1;
    (* src = "src/sreg.spade:27,19" *)
    logic val_n2;
    (* src = "src/sreg.spade:29,19" *)
    logic val_n3;
    (* src = "src/sreg.spade:31,19" *)
    logic val_n4;
    (* src = "src/sreg.spade:33,19" *)
    logic val_n5;
    (* src = "src/sreg.spade:35,19" *)
    logic val_n6;
    (* src = "src/sreg.spade:37,19" *)
    logic val_n7;
    (* src = "src/sreg.spade:39,19" *)
    logic val_n8;
    (* src = "src/sreg.spade:41,19" *)
    logic val_n9;
    (* src = "src/sreg.spade:43,19" *)
    logic val_n10;
    (* src = "src/sreg.spade:45,19" *)
    logic val_n11;
    (* src = "src/sreg.spade:47,19" *)
    logic val_n12;
    (* src = "src/sreg.spade:49,19" *)
    logic val_n13;
    (* src = "src/sreg.spade:51,19" *)
    logic val_n14;
    (* src = "src/sreg.spade:53,19" *)
    logic val_n15;
    (* src = "src/sreg.spade:55,19" *)
    logic val_n16;
    (* src = "src/sreg.spade:57,19" *)
    logic val_n17;
    (* src = "src/sreg.spade:59,19" *)
    logic val_n18;
    (* src = "src/sreg.spade:61,19" *)
    logic val_n19;
    (* src = "src/sreg.spade:63,19" *)
    logic val_n20;
    (* src = "src/sreg.spade:65,19" *)
    logic val_n21;
    (* src = "src/sreg.spade:67,19" *)
    logic val_n22;
    (* src = "src/sreg.spade:69,19" *)
    logic val_n23;
    (* src = "src/sreg.spade:71,19" *)
    logic val_n24;
    (* src = "src/sreg.spade:73,19" *)
    logic val_n25;
    (* src = "src/sreg.spade:75,19" *)
    logic val_n26;
    (* src = "src/sreg.spade:77,19" *)
    logic val_n27;
    (* src = "src/sreg.spade:79,19" *)
    logic val_n28;
    (* src = "src/sreg.spade:81,19" *)
    logic val_n29;
    (* src = "src/sreg.spade:83,19" *)
    logic val_n30;
    (* src = "src/sreg.spade:85,19" *)
    logic val_n31;
    (* src = "src/sreg.spade:87,19" *)
    logic val_n32;
    (* src = "src/sreg.spade:89,19" *)
    logic val_n33;
    (* src = "src/sreg.spade:91,19" *)
    logic val_n34;
    (* src = "src/sreg.spade:93,19" *)
    logic val_n35;
    (* src = "src/sreg.spade:95,19" *)
    logic val_n36;
    (* src = "src/sreg.spade:97,19" *)
    logic val_n37;
    (* src = "src/sreg.spade:99,19" *)
    logic val_n38;
    (* src = "src/sreg.spade:101,19" *)
    logic val_n39;
    (* src = "src/sreg.spade:103,19" *)
    logic val_n40;
    (* src = "src/sreg.spade:105,19" *)
    logic val_n41;
    (* src = "src/sreg.spade:107,19" *)
    logic val_n42;
    (* src = "src/sreg.spade:109,19" *)
    logic val_n43;
    (* src = "src/sreg.spade:111,19" *)
    logic val_n44;
    (* src = "src/sreg.spade:113,19" *)
    logic val_n45;
    (* src = "src/sreg.spade:115,19" *)
    logic val_n46;
    (* src = "src/sreg.spade:117,19" *)
    logic val_n47;
    (* src = "src/sreg.spade:119,19" *)
    logic val_n48;
    (* src = "src/sreg.spade:121,19" *)
    logic val_n49;
    always @(posedge \clk ) begin
        \s1_val  <= \val ;
    end
    always @(posedge \clk ) begin
        \s2_val  <= \s1_val ;
    end
    always @(posedge \clk ) begin
        \s3_val  <= \s2_val ;
    end
    always @(posedge \clk ) begin
        \s4_val  <= \s3_val ;
    end
    always @(posedge \clk ) begin
        \s5_val  <= \s4_val ;
    end
    always @(posedge \clk ) begin
        s5_val_n1 <= val_n1;
    end
    always @(posedge \clk ) begin
        \s6_val  <= \s5_val ;
    end
    always @(posedge \clk ) begin
        s6_val_n1 <= s5_val_n1;
    end
    always @(posedge \clk ) begin
        \s7_val  <= \s6_val ;
    end
    always @(posedge \clk ) begin
        s7_val_n1 <= s6_val_n1;
    end
    always @(posedge \clk ) begin
        s7_val_n2 <= val_n2;
    end
    always @(posedge \clk ) begin
        \s8_val  <= \s7_val ;
    end
    always @(posedge \clk ) begin
        s8_val_n1 <= s7_val_n1;
    end
    always @(posedge \clk ) begin
        s8_val_n2 <= s7_val_n2;
    end
    always @(posedge \clk ) begin
        \s9_val  <= \s8_val ;
    end
    always @(posedge \clk ) begin
        s9_val_n1 <= s8_val_n1;
    end
    always @(posedge \clk ) begin
        s9_val_n2 <= s8_val_n2;
    end
    always @(posedge \clk ) begin
        s9_val_n3 <= val_n3;
    end
    always @(posedge \clk ) begin
        \s10_val  <= \s9_val ;
    end
    always @(posedge \clk ) begin
        s10_val_n1 <= s9_val_n1;
    end
    always @(posedge \clk ) begin
        s10_val_n2 <= s9_val_n2;
    end
    always @(posedge \clk ) begin
        s10_val_n3 <= s9_val_n3;
    end
    always @(posedge \clk ) begin
        \s11_val  <= \s10_val ;
    end
    always @(posedge \clk ) begin
        s11_val_n1 <= s10_val_n1;
    end
    always @(posedge \clk ) begin
        s11_val_n2 <= s10_val_n2;
    end
    always @(posedge \clk ) begin
        s11_val_n3 <= s10_val_n3;
    end
    always @(posedge \clk ) begin
        s11_val_n4 <= val_n4;
    end
    always @(posedge \clk ) begin
        \s12_val  <= \s11_val ;
    end
    always @(posedge \clk ) begin
        s12_val_n1 <= s11_val_n1;
    end
    always @(posedge \clk ) begin
        s12_val_n2 <= s11_val_n2;
    end
    always @(posedge \clk ) begin
        s12_val_n3 <= s11_val_n3;
    end
    always @(posedge \clk ) begin
        s12_val_n4 <= s11_val_n4;
    end
    always @(posedge \clk ) begin
        \s13_val  <= \s12_val ;
    end
    always @(posedge \clk ) begin
        s13_val_n1 <= s12_val_n1;
    end
    always @(posedge \clk ) begin
        s13_val_n2 <= s12_val_n2;
    end
    always @(posedge \clk ) begin
        s13_val_n3 <= s12_val_n3;
    end
    always @(posedge \clk ) begin
        s13_val_n4 <= s12_val_n4;
    end
    always @(posedge \clk ) begin
        s13_val_n5 <= val_n5;
    end
    always @(posedge \clk ) begin
        \s14_val  <= \s13_val ;
    end
    always @(posedge \clk ) begin
        s14_val_n1 <= s13_val_n1;
    end
    always @(posedge \clk ) begin
        s14_val_n2 <= s13_val_n2;
    end
    always @(posedge \clk ) begin
        s14_val_n3 <= s13_val_n3;
    end
    always @(posedge \clk ) begin
        s14_val_n4 <= s13_val_n4;
    end
    always @(posedge \clk ) begin
        s14_val_n5 <= s13_val_n5;
    end
    always @(posedge \clk ) begin
        \s15_val  <= \s14_val ;
    end
    always @(posedge \clk ) begin
        s15_val_n1 <= s14_val_n1;
    end
    always @(posedge \clk ) begin
        s15_val_n2 <= s14_val_n2;
    end
    always @(posedge \clk ) begin
        s15_val_n3 <= s14_val_n3;
    end
    always @(posedge \clk ) begin
        s15_val_n4 <= s14_val_n4;
    end
    always @(posedge \clk ) begin
        s15_val_n5 <= s14_val_n5;
    end
    always @(posedge \clk ) begin
        s15_val_n6 <= val_n6;
    end
    always @(posedge \clk ) begin
        \s16_val  <= \s15_val ;
    end
    always @(posedge \clk ) begin
        s16_val_n1 <= s15_val_n1;
    end
    always @(posedge \clk ) begin
        s16_val_n2 <= s15_val_n2;
    end
    always @(posedge \clk ) begin
        s16_val_n3 <= s15_val_n3;
    end
    always @(posedge \clk ) begin
        s16_val_n4 <= s15_val_n4;
    end
    always @(posedge \clk ) begin
        s16_val_n5 <= s15_val_n5;
    end
    always @(posedge \clk ) begin
        s16_val_n6 <= s15_val_n6;
    end
    always @(posedge \clk ) begin
        \s17_val  <= \s16_val ;
    end
    always @(posedge \clk ) begin
        s17_val_n1 <= s16_val_n1;
    end
    always @(posedge \clk ) begin
        s17_val_n2 <= s16_val_n2;
    end
    always @(posedge \clk ) begin
        s17_val_n3 <= s16_val_n3;
    end
    always @(posedge \clk ) begin
        s17_val_n4 <= s16_val_n4;
    end
    always @(posedge \clk ) begin
        s17_val_n5 <= s16_val_n5;
    end
    always @(posedge \clk ) begin
        s17_val_n6 <= s16_val_n6;
    end
    always @(posedge \clk ) begin
        s17_val_n7 <= val_n7;
    end
    always @(posedge \clk ) begin
        \s18_val  <= \s17_val ;
    end
    always @(posedge \clk ) begin
        s18_val_n1 <= s17_val_n1;
    end
    always @(posedge \clk ) begin
        s18_val_n2 <= s17_val_n2;
    end
    always @(posedge \clk ) begin
        s18_val_n3 <= s17_val_n3;
    end
    always @(posedge \clk ) begin
        s18_val_n4 <= s17_val_n4;
    end
    always @(posedge \clk ) begin
        s18_val_n5 <= s17_val_n5;
    end
    always @(posedge \clk ) begin
        s18_val_n6 <= s17_val_n6;
    end
    always @(posedge \clk ) begin
        s18_val_n7 <= s17_val_n7;
    end
    always @(posedge \clk ) begin
        \s19_val  <= \s18_val ;
    end
    always @(posedge \clk ) begin
        s19_val_n1 <= s18_val_n1;
    end
    always @(posedge \clk ) begin
        s19_val_n2 <= s18_val_n2;
    end
    always @(posedge \clk ) begin
        s19_val_n3 <= s18_val_n3;
    end
    always @(posedge \clk ) begin
        s19_val_n4 <= s18_val_n4;
    end
    always @(posedge \clk ) begin
        s19_val_n5 <= s18_val_n5;
    end
    always @(posedge \clk ) begin
        s19_val_n6 <= s18_val_n6;
    end
    always @(posedge \clk ) begin
        s19_val_n7 <= s18_val_n7;
    end
    always @(posedge \clk ) begin
        s19_val_n8 <= val_n8;
    end
    always @(posedge \clk ) begin
        \s20_val  <= \s19_val ;
    end
    always @(posedge \clk ) begin
        s20_val_n1 <= s19_val_n1;
    end
    always @(posedge \clk ) begin
        s20_val_n2 <= s19_val_n2;
    end
    always @(posedge \clk ) begin
        s20_val_n3 <= s19_val_n3;
    end
    always @(posedge \clk ) begin
        s20_val_n4 <= s19_val_n4;
    end
    always @(posedge \clk ) begin
        s20_val_n5 <= s19_val_n5;
    end
    always @(posedge \clk ) begin
        s20_val_n6 <= s19_val_n6;
    end
    always @(posedge \clk ) begin
        s20_val_n7 <= s19_val_n7;
    end
    always @(posedge \clk ) begin
        s20_val_n8 <= s19_val_n8;
    end
    always @(posedge \clk ) begin
        \s21_val  <= \s20_val ;
    end
    always @(posedge \clk ) begin
        s21_val_n1 <= s20_val_n1;
    end
    always @(posedge \clk ) begin
        s21_val_n2 <= s20_val_n2;
    end
    always @(posedge \clk ) begin
        s21_val_n3 <= s20_val_n3;
    end
    always @(posedge \clk ) begin
        s21_val_n4 <= s20_val_n4;
    end
    always @(posedge \clk ) begin
        s21_val_n5 <= s20_val_n5;
    end
    always @(posedge \clk ) begin
        s21_val_n6 <= s20_val_n6;
    end
    always @(posedge \clk ) begin
        s21_val_n7 <= s20_val_n7;
    end
    always @(posedge \clk ) begin
        s21_val_n8 <= s20_val_n8;
    end
    always @(posedge \clk ) begin
        s21_val_n9 <= val_n9;
    end
    always @(posedge \clk ) begin
        \s22_val  <= \s21_val ;
    end
    always @(posedge \clk ) begin
        s22_val_n1 <= s21_val_n1;
    end
    always @(posedge \clk ) begin
        s22_val_n2 <= s21_val_n2;
    end
    always @(posedge \clk ) begin
        s22_val_n3 <= s21_val_n3;
    end
    always @(posedge \clk ) begin
        s22_val_n4 <= s21_val_n4;
    end
    always @(posedge \clk ) begin
        s22_val_n5 <= s21_val_n5;
    end
    always @(posedge \clk ) begin
        s22_val_n6 <= s21_val_n6;
    end
    always @(posedge \clk ) begin
        s22_val_n7 <= s21_val_n7;
    end
    always @(posedge \clk ) begin
        s22_val_n8 <= s21_val_n8;
    end
    always @(posedge \clk ) begin
        s22_val_n9 <= s21_val_n9;
    end
    always @(posedge \clk ) begin
        \s23_val  <= \s22_val ;
    end
    always @(posedge \clk ) begin
        s23_val_n1 <= s22_val_n1;
    end
    always @(posedge \clk ) begin
        s23_val_n2 <= s22_val_n2;
    end
    always @(posedge \clk ) begin
        s23_val_n3 <= s22_val_n3;
    end
    always @(posedge \clk ) begin
        s23_val_n4 <= s22_val_n4;
    end
    always @(posedge \clk ) begin
        s23_val_n5 <= s22_val_n5;
    end
    always @(posedge \clk ) begin
        s23_val_n6 <= s22_val_n6;
    end
    always @(posedge \clk ) begin
        s23_val_n7 <= s22_val_n7;
    end
    always @(posedge \clk ) begin
        s23_val_n8 <= s22_val_n8;
    end
    always @(posedge \clk ) begin
        s23_val_n9 <= s22_val_n9;
    end
    always @(posedge \clk ) begin
        s23_val_n10 <= val_n10;
    end
    always @(posedge \clk ) begin
        \s24_val  <= \s23_val ;
    end
    always @(posedge \clk ) begin
        s24_val_n1 <= s23_val_n1;
    end
    always @(posedge \clk ) begin
        s24_val_n2 <= s23_val_n2;
    end
    always @(posedge \clk ) begin
        s24_val_n3 <= s23_val_n3;
    end
    always @(posedge \clk ) begin
        s24_val_n4 <= s23_val_n4;
    end
    always @(posedge \clk ) begin
        s24_val_n5 <= s23_val_n5;
    end
    always @(posedge \clk ) begin
        s24_val_n6 <= s23_val_n6;
    end
    always @(posedge \clk ) begin
        s24_val_n7 <= s23_val_n7;
    end
    always @(posedge \clk ) begin
        s24_val_n8 <= s23_val_n8;
    end
    always @(posedge \clk ) begin
        s24_val_n9 <= s23_val_n9;
    end
    always @(posedge \clk ) begin
        s24_val_n10 <= s23_val_n10;
    end
    always @(posedge \clk ) begin
        \s25_val  <= \s24_val ;
    end
    always @(posedge \clk ) begin
        s25_val_n1 <= s24_val_n1;
    end
    always @(posedge \clk ) begin
        s25_val_n2 <= s24_val_n2;
    end
    always @(posedge \clk ) begin
        s25_val_n3 <= s24_val_n3;
    end
    always @(posedge \clk ) begin
        s25_val_n4 <= s24_val_n4;
    end
    always @(posedge \clk ) begin
        s25_val_n5 <= s24_val_n5;
    end
    always @(posedge \clk ) begin
        s25_val_n6 <= s24_val_n6;
    end
    always @(posedge \clk ) begin
        s25_val_n7 <= s24_val_n7;
    end
    always @(posedge \clk ) begin
        s25_val_n8 <= s24_val_n8;
    end
    always @(posedge \clk ) begin
        s25_val_n9 <= s24_val_n9;
    end
    always @(posedge \clk ) begin
        s25_val_n10 <= s24_val_n10;
    end
    always @(posedge \clk ) begin
        s25_val_n11 <= val_n11;
    end
    always @(posedge \clk ) begin
        \s26_val  <= \s25_val ;
    end
    always @(posedge \clk ) begin
        s26_val_n1 <= s25_val_n1;
    end
    always @(posedge \clk ) begin
        s26_val_n2 <= s25_val_n2;
    end
    always @(posedge \clk ) begin
        s26_val_n3 <= s25_val_n3;
    end
    always @(posedge \clk ) begin
        s26_val_n4 <= s25_val_n4;
    end
    always @(posedge \clk ) begin
        s26_val_n5 <= s25_val_n5;
    end
    always @(posedge \clk ) begin
        s26_val_n6 <= s25_val_n6;
    end
    always @(posedge \clk ) begin
        s26_val_n7 <= s25_val_n7;
    end
    always @(posedge \clk ) begin
        s26_val_n8 <= s25_val_n8;
    end
    always @(posedge \clk ) begin
        s26_val_n9 <= s25_val_n9;
    end
    always @(posedge \clk ) begin
        s26_val_n10 <= s25_val_n10;
    end
    always @(posedge \clk ) begin
        s26_val_n11 <= s25_val_n11;
    end
    always @(posedge \clk ) begin
        \s27_val  <= \s26_val ;
    end
    always @(posedge \clk ) begin
        s27_val_n1 <= s26_val_n1;
    end
    always @(posedge \clk ) begin
        s27_val_n2 <= s26_val_n2;
    end
    always @(posedge \clk ) begin
        s27_val_n3 <= s26_val_n3;
    end
    always @(posedge \clk ) begin
        s27_val_n4 <= s26_val_n4;
    end
    always @(posedge \clk ) begin
        s27_val_n5 <= s26_val_n5;
    end
    always @(posedge \clk ) begin
        s27_val_n6 <= s26_val_n6;
    end
    always @(posedge \clk ) begin
        s27_val_n7 <= s26_val_n7;
    end
    always @(posedge \clk ) begin
        s27_val_n8 <= s26_val_n8;
    end
    always @(posedge \clk ) begin
        s27_val_n9 <= s26_val_n9;
    end
    always @(posedge \clk ) begin
        s27_val_n10 <= s26_val_n10;
    end
    always @(posedge \clk ) begin
        s27_val_n11 <= s26_val_n11;
    end
    always @(posedge \clk ) begin
        s27_val_n12 <= val_n12;
    end
    always @(posedge \clk ) begin
        \s28_val  <= \s27_val ;
    end
    always @(posedge \clk ) begin
        s28_val_n1 <= s27_val_n1;
    end
    always @(posedge \clk ) begin
        s28_val_n2 <= s27_val_n2;
    end
    always @(posedge \clk ) begin
        s28_val_n3 <= s27_val_n3;
    end
    always @(posedge \clk ) begin
        s28_val_n4 <= s27_val_n4;
    end
    always @(posedge \clk ) begin
        s28_val_n5 <= s27_val_n5;
    end
    always @(posedge \clk ) begin
        s28_val_n6 <= s27_val_n6;
    end
    always @(posedge \clk ) begin
        s28_val_n7 <= s27_val_n7;
    end
    always @(posedge \clk ) begin
        s28_val_n8 <= s27_val_n8;
    end
    always @(posedge \clk ) begin
        s28_val_n9 <= s27_val_n9;
    end
    always @(posedge \clk ) begin
        s28_val_n10 <= s27_val_n10;
    end
    always @(posedge \clk ) begin
        s28_val_n11 <= s27_val_n11;
    end
    always @(posedge \clk ) begin
        s28_val_n12 <= s27_val_n12;
    end
    always @(posedge \clk ) begin
        \s29_val  <= \s28_val ;
    end
    always @(posedge \clk ) begin
        s29_val_n1 <= s28_val_n1;
    end
    always @(posedge \clk ) begin
        s29_val_n2 <= s28_val_n2;
    end
    always @(posedge \clk ) begin
        s29_val_n3 <= s28_val_n3;
    end
    always @(posedge \clk ) begin
        s29_val_n4 <= s28_val_n4;
    end
    always @(posedge \clk ) begin
        s29_val_n5 <= s28_val_n5;
    end
    always @(posedge \clk ) begin
        s29_val_n6 <= s28_val_n6;
    end
    always @(posedge \clk ) begin
        s29_val_n7 <= s28_val_n7;
    end
    always @(posedge \clk ) begin
        s29_val_n8 <= s28_val_n8;
    end
    always @(posedge \clk ) begin
        s29_val_n9 <= s28_val_n9;
    end
    always @(posedge \clk ) begin
        s29_val_n10 <= s28_val_n10;
    end
    always @(posedge \clk ) begin
        s29_val_n11 <= s28_val_n11;
    end
    always @(posedge \clk ) begin
        s29_val_n12 <= s28_val_n12;
    end
    always @(posedge \clk ) begin
        s29_val_n13 <= val_n13;
    end
    always @(posedge \clk ) begin
        \s30_val  <= \s29_val ;
    end
    always @(posedge \clk ) begin
        s30_val_n1 <= s29_val_n1;
    end
    always @(posedge \clk ) begin
        s30_val_n2 <= s29_val_n2;
    end
    always @(posedge \clk ) begin
        s30_val_n3 <= s29_val_n3;
    end
    always @(posedge \clk ) begin
        s30_val_n4 <= s29_val_n4;
    end
    always @(posedge \clk ) begin
        s30_val_n5 <= s29_val_n5;
    end
    always @(posedge \clk ) begin
        s30_val_n6 <= s29_val_n6;
    end
    always @(posedge \clk ) begin
        s30_val_n7 <= s29_val_n7;
    end
    always @(posedge \clk ) begin
        s30_val_n8 <= s29_val_n8;
    end
    always @(posedge \clk ) begin
        s30_val_n9 <= s29_val_n9;
    end
    always @(posedge \clk ) begin
        s30_val_n10 <= s29_val_n10;
    end
    always @(posedge \clk ) begin
        s30_val_n11 <= s29_val_n11;
    end
    always @(posedge \clk ) begin
        s30_val_n12 <= s29_val_n12;
    end
    always @(posedge \clk ) begin
        s30_val_n13 <= s29_val_n13;
    end
    always @(posedge \clk ) begin
        \s31_val  <= \s30_val ;
    end
    always @(posedge \clk ) begin
        s31_val_n1 <= s30_val_n1;
    end
    always @(posedge \clk ) begin
        s31_val_n2 <= s30_val_n2;
    end
    always @(posedge \clk ) begin
        s31_val_n3 <= s30_val_n3;
    end
    always @(posedge \clk ) begin
        s31_val_n4 <= s30_val_n4;
    end
    always @(posedge \clk ) begin
        s31_val_n5 <= s30_val_n5;
    end
    always @(posedge \clk ) begin
        s31_val_n6 <= s30_val_n6;
    end
    always @(posedge \clk ) begin
        s31_val_n7 <= s30_val_n7;
    end
    always @(posedge \clk ) begin
        s31_val_n8 <= s30_val_n8;
    end
    always @(posedge \clk ) begin
        s31_val_n9 <= s30_val_n9;
    end
    always @(posedge \clk ) begin
        s31_val_n10 <= s30_val_n10;
    end
    always @(posedge \clk ) begin
        s31_val_n11 <= s30_val_n11;
    end
    always @(posedge \clk ) begin
        s31_val_n12 <= s30_val_n12;
    end
    always @(posedge \clk ) begin
        s31_val_n13 <= s30_val_n13;
    end
    always @(posedge \clk ) begin
        s31_val_n14 <= val_n14;
    end
    always @(posedge \clk ) begin
        \s32_val  <= \s31_val ;
    end
    always @(posedge \clk ) begin
        s32_val_n1 <= s31_val_n1;
    end
    always @(posedge \clk ) begin
        s32_val_n2 <= s31_val_n2;
    end
    always @(posedge \clk ) begin
        s32_val_n3 <= s31_val_n3;
    end
    always @(posedge \clk ) begin
        s32_val_n4 <= s31_val_n4;
    end
    always @(posedge \clk ) begin
        s32_val_n5 <= s31_val_n5;
    end
    always @(posedge \clk ) begin
        s32_val_n6 <= s31_val_n6;
    end
    always @(posedge \clk ) begin
        s32_val_n7 <= s31_val_n7;
    end
    always @(posedge \clk ) begin
        s32_val_n8 <= s31_val_n8;
    end
    always @(posedge \clk ) begin
        s32_val_n9 <= s31_val_n9;
    end
    always @(posedge \clk ) begin
        s32_val_n10 <= s31_val_n10;
    end
    always @(posedge \clk ) begin
        s32_val_n11 <= s31_val_n11;
    end
    always @(posedge \clk ) begin
        s32_val_n12 <= s31_val_n12;
    end
    always @(posedge \clk ) begin
        s32_val_n13 <= s31_val_n13;
    end
    always @(posedge \clk ) begin
        s32_val_n14 <= s31_val_n14;
    end
    always @(posedge \clk ) begin
        \s33_val  <= \s32_val ;
    end
    always @(posedge \clk ) begin
        s33_val_n1 <= s32_val_n1;
    end
    always @(posedge \clk ) begin
        s33_val_n2 <= s32_val_n2;
    end
    always @(posedge \clk ) begin
        s33_val_n3 <= s32_val_n3;
    end
    always @(posedge \clk ) begin
        s33_val_n4 <= s32_val_n4;
    end
    always @(posedge \clk ) begin
        s33_val_n5 <= s32_val_n5;
    end
    always @(posedge \clk ) begin
        s33_val_n6 <= s32_val_n6;
    end
    always @(posedge \clk ) begin
        s33_val_n7 <= s32_val_n7;
    end
    always @(posedge \clk ) begin
        s33_val_n8 <= s32_val_n8;
    end
    always @(posedge \clk ) begin
        s33_val_n9 <= s32_val_n9;
    end
    always @(posedge \clk ) begin
        s33_val_n10 <= s32_val_n10;
    end
    always @(posedge \clk ) begin
        s33_val_n11 <= s32_val_n11;
    end
    always @(posedge \clk ) begin
        s33_val_n12 <= s32_val_n12;
    end
    always @(posedge \clk ) begin
        s33_val_n13 <= s32_val_n13;
    end
    always @(posedge \clk ) begin
        s33_val_n14 <= s32_val_n14;
    end
    always @(posedge \clk ) begin
        s33_val_n15 <= val_n15;
    end
    always @(posedge \clk ) begin
        \s34_val  <= \s33_val ;
    end
    always @(posedge \clk ) begin
        s34_val_n1 <= s33_val_n1;
    end
    always @(posedge \clk ) begin
        s34_val_n2 <= s33_val_n2;
    end
    always @(posedge \clk ) begin
        s34_val_n3 <= s33_val_n3;
    end
    always @(posedge \clk ) begin
        s34_val_n4 <= s33_val_n4;
    end
    always @(posedge \clk ) begin
        s34_val_n5 <= s33_val_n5;
    end
    always @(posedge \clk ) begin
        s34_val_n6 <= s33_val_n6;
    end
    always @(posedge \clk ) begin
        s34_val_n7 <= s33_val_n7;
    end
    always @(posedge \clk ) begin
        s34_val_n8 <= s33_val_n8;
    end
    always @(posedge \clk ) begin
        s34_val_n9 <= s33_val_n9;
    end
    always @(posedge \clk ) begin
        s34_val_n10 <= s33_val_n10;
    end
    always @(posedge \clk ) begin
        s34_val_n11 <= s33_val_n11;
    end
    always @(posedge \clk ) begin
        s34_val_n12 <= s33_val_n12;
    end
    always @(posedge \clk ) begin
        s34_val_n13 <= s33_val_n13;
    end
    always @(posedge \clk ) begin
        s34_val_n14 <= s33_val_n14;
    end
    always @(posedge \clk ) begin
        s34_val_n15 <= s33_val_n15;
    end
    always @(posedge \clk ) begin
        \s35_val  <= \s34_val ;
    end
    always @(posedge \clk ) begin
        s35_val_n1 <= s34_val_n1;
    end
    always @(posedge \clk ) begin
        s35_val_n2 <= s34_val_n2;
    end
    always @(posedge \clk ) begin
        s35_val_n3 <= s34_val_n3;
    end
    always @(posedge \clk ) begin
        s35_val_n4 <= s34_val_n4;
    end
    always @(posedge \clk ) begin
        s35_val_n5 <= s34_val_n5;
    end
    always @(posedge \clk ) begin
        s35_val_n6 <= s34_val_n6;
    end
    always @(posedge \clk ) begin
        s35_val_n7 <= s34_val_n7;
    end
    always @(posedge \clk ) begin
        s35_val_n8 <= s34_val_n8;
    end
    always @(posedge \clk ) begin
        s35_val_n9 <= s34_val_n9;
    end
    always @(posedge \clk ) begin
        s35_val_n10 <= s34_val_n10;
    end
    always @(posedge \clk ) begin
        s35_val_n11 <= s34_val_n11;
    end
    always @(posedge \clk ) begin
        s35_val_n12 <= s34_val_n12;
    end
    always @(posedge \clk ) begin
        s35_val_n13 <= s34_val_n13;
    end
    always @(posedge \clk ) begin
        s35_val_n14 <= s34_val_n14;
    end
    always @(posedge \clk ) begin
        s35_val_n15 <= s34_val_n15;
    end
    always @(posedge \clk ) begin
        s35_val_n16 <= val_n16;
    end
    always @(posedge \clk ) begin
        \s36_val  <= \s35_val ;
    end
    always @(posedge \clk ) begin
        s36_val_n1 <= s35_val_n1;
    end
    always @(posedge \clk ) begin
        s36_val_n2 <= s35_val_n2;
    end
    always @(posedge \clk ) begin
        s36_val_n3 <= s35_val_n3;
    end
    always @(posedge \clk ) begin
        s36_val_n4 <= s35_val_n4;
    end
    always @(posedge \clk ) begin
        s36_val_n5 <= s35_val_n5;
    end
    always @(posedge \clk ) begin
        s36_val_n6 <= s35_val_n6;
    end
    always @(posedge \clk ) begin
        s36_val_n7 <= s35_val_n7;
    end
    always @(posedge \clk ) begin
        s36_val_n8 <= s35_val_n8;
    end
    always @(posedge \clk ) begin
        s36_val_n9 <= s35_val_n9;
    end
    always @(posedge \clk ) begin
        s36_val_n10 <= s35_val_n10;
    end
    always @(posedge \clk ) begin
        s36_val_n11 <= s35_val_n11;
    end
    always @(posedge \clk ) begin
        s36_val_n12 <= s35_val_n12;
    end
    always @(posedge \clk ) begin
        s36_val_n13 <= s35_val_n13;
    end
    always @(posedge \clk ) begin
        s36_val_n14 <= s35_val_n14;
    end
    always @(posedge \clk ) begin
        s36_val_n15 <= s35_val_n15;
    end
    always @(posedge \clk ) begin
        s36_val_n16 <= s35_val_n16;
    end
    always @(posedge \clk ) begin
        \s37_val  <= \s36_val ;
    end
    always @(posedge \clk ) begin
        s37_val_n1 <= s36_val_n1;
    end
    always @(posedge \clk ) begin
        s37_val_n2 <= s36_val_n2;
    end
    always @(posedge \clk ) begin
        s37_val_n3 <= s36_val_n3;
    end
    always @(posedge \clk ) begin
        s37_val_n4 <= s36_val_n4;
    end
    always @(posedge \clk ) begin
        s37_val_n5 <= s36_val_n5;
    end
    always @(posedge \clk ) begin
        s37_val_n6 <= s36_val_n6;
    end
    always @(posedge \clk ) begin
        s37_val_n7 <= s36_val_n7;
    end
    always @(posedge \clk ) begin
        s37_val_n8 <= s36_val_n8;
    end
    always @(posedge \clk ) begin
        s37_val_n9 <= s36_val_n9;
    end
    always @(posedge \clk ) begin
        s37_val_n10 <= s36_val_n10;
    end
    always @(posedge \clk ) begin
        s37_val_n11 <= s36_val_n11;
    end
    always @(posedge \clk ) begin
        s37_val_n12 <= s36_val_n12;
    end
    always @(posedge \clk ) begin
        s37_val_n13 <= s36_val_n13;
    end
    always @(posedge \clk ) begin
        s37_val_n14 <= s36_val_n14;
    end
    always @(posedge \clk ) begin
        s37_val_n15 <= s36_val_n15;
    end
    always @(posedge \clk ) begin
        s37_val_n16 <= s36_val_n16;
    end
    always @(posedge \clk ) begin
        s37_val_n17 <= val_n17;
    end
    always @(posedge \clk ) begin
        \s38_val  <= \s37_val ;
    end
    always @(posedge \clk ) begin
        s38_val_n1 <= s37_val_n1;
    end
    always @(posedge \clk ) begin
        s38_val_n2 <= s37_val_n2;
    end
    always @(posedge \clk ) begin
        s38_val_n3 <= s37_val_n3;
    end
    always @(posedge \clk ) begin
        s38_val_n4 <= s37_val_n4;
    end
    always @(posedge \clk ) begin
        s38_val_n5 <= s37_val_n5;
    end
    always @(posedge \clk ) begin
        s38_val_n6 <= s37_val_n6;
    end
    always @(posedge \clk ) begin
        s38_val_n7 <= s37_val_n7;
    end
    always @(posedge \clk ) begin
        s38_val_n8 <= s37_val_n8;
    end
    always @(posedge \clk ) begin
        s38_val_n9 <= s37_val_n9;
    end
    always @(posedge \clk ) begin
        s38_val_n10 <= s37_val_n10;
    end
    always @(posedge \clk ) begin
        s38_val_n11 <= s37_val_n11;
    end
    always @(posedge \clk ) begin
        s38_val_n12 <= s37_val_n12;
    end
    always @(posedge \clk ) begin
        s38_val_n13 <= s37_val_n13;
    end
    always @(posedge \clk ) begin
        s38_val_n14 <= s37_val_n14;
    end
    always @(posedge \clk ) begin
        s38_val_n15 <= s37_val_n15;
    end
    always @(posedge \clk ) begin
        s38_val_n16 <= s37_val_n16;
    end
    always @(posedge \clk ) begin
        s38_val_n17 <= s37_val_n17;
    end
    always @(posedge \clk ) begin
        \s39_val  <= \s38_val ;
    end
    always @(posedge \clk ) begin
        s39_val_n1 <= s38_val_n1;
    end
    always @(posedge \clk ) begin
        s39_val_n2 <= s38_val_n2;
    end
    always @(posedge \clk ) begin
        s39_val_n3 <= s38_val_n3;
    end
    always @(posedge \clk ) begin
        s39_val_n4 <= s38_val_n4;
    end
    always @(posedge \clk ) begin
        s39_val_n5 <= s38_val_n5;
    end
    always @(posedge \clk ) begin
        s39_val_n6 <= s38_val_n6;
    end
    always @(posedge \clk ) begin
        s39_val_n7 <= s38_val_n7;
    end
    always @(posedge \clk ) begin
        s39_val_n8 <= s38_val_n8;
    end
    always @(posedge \clk ) begin
        s39_val_n9 <= s38_val_n9;
    end
    always @(posedge \clk ) begin
        s39_val_n10 <= s38_val_n10;
    end
    always @(posedge \clk ) begin
        s39_val_n11 <= s38_val_n11;
    end
    always @(posedge \clk ) begin
        s39_val_n12 <= s38_val_n12;
    end
    always @(posedge \clk ) begin
        s39_val_n13 <= s38_val_n13;
    end
    always @(posedge \clk ) begin
        s39_val_n14 <= s38_val_n14;
    end
    always @(posedge \clk ) begin
        s39_val_n15 <= s38_val_n15;
    end
    always @(posedge \clk ) begin
        s39_val_n16 <= s38_val_n16;
    end
    always @(posedge \clk ) begin
        s39_val_n17 <= s38_val_n17;
    end
    always @(posedge \clk ) begin
        s39_val_n18 <= val_n18;
    end
    always @(posedge \clk ) begin
        \s40_val  <= \s39_val ;
    end
    always @(posedge \clk ) begin
        s40_val_n1 <= s39_val_n1;
    end
    always @(posedge \clk ) begin
        s40_val_n2 <= s39_val_n2;
    end
    always @(posedge \clk ) begin
        s40_val_n3 <= s39_val_n3;
    end
    always @(posedge \clk ) begin
        s40_val_n4 <= s39_val_n4;
    end
    always @(posedge \clk ) begin
        s40_val_n5 <= s39_val_n5;
    end
    always @(posedge \clk ) begin
        s40_val_n6 <= s39_val_n6;
    end
    always @(posedge \clk ) begin
        s40_val_n7 <= s39_val_n7;
    end
    always @(posedge \clk ) begin
        s40_val_n8 <= s39_val_n8;
    end
    always @(posedge \clk ) begin
        s40_val_n9 <= s39_val_n9;
    end
    always @(posedge \clk ) begin
        s40_val_n10 <= s39_val_n10;
    end
    always @(posedge \clk ) begin
        s40_val_n11 <= s39_val_n11;
    end
    always @(posedge \clk ) begin
        s40_val_n12 <= s39_val_n12;
    end
    always @(posedge \clk ) begin
        s40_val_n13 <= s39_val_n13;
    end
    always @(posedge \clk ) begin
        s40_val_n14 <= s39_val_n14;
    end
    always @(posedge \clk ) begin
        s40_val_n15 <= s39_val_n15;
    end
    always @(posedge \clk ) begin
        s40_val_n16 <= s39_val_n16;
    end
    always @(posedge \clk ) begin
        s40_val_n17 <= s39_val_n17;
    end
    always @(posedge \clk ) begin
        s40_val_n18 <= s39_val_n18;
    end
    always @(posedge \clk ) begin
        \s41_val  <= \s40_val ;
    end
    always @(posedge \clk ) begin
        s41_val_n1 <= s40_val_n1;
    end
    always @(posedge \clk ) begin
        s41_val_n2 <= s40_val_n2;
    end
    always @(posedge \clk ) begin
        s41_val_n3 <= s40_val_n3;
    end
    always @(posedge \clk ) begin
        s41_val_n4 <= s40_val_n4;
    end
    always @(posedge \clk ) begin
        s41_val_n5 <= s40_val_n5;
    end
    always @(posedge \clk ) begin
        s41_val_n6 <= s40_val_n6;
    end
    always @(posedge \clk ) begin
        s41_val_n7 <= s40_val_n7;
    end
    always @(posedge \clk ) begin
        s41_val_n8 <= s40_val_n8;
    end
    always @(posedge \clk ) begin
        s41_val_n9 <= s40_val_n9;
    end
    always @(posedge \clk ) begin
        s41_val_n10 <= s40_val_n10;
    end
    always @(posedge \clk ) begin
        s41_val_n11 <= s40_val_n11;
    end
    always @(posedge \clk ) begin
        s41_val_n12 <= s40_val_n12;
    end
    always @(posedge \clk ) begin
        s41_val_n13 <= s40_val_n13;
    end
    always @(posedge \clk ) begin
        s41_val_n14 <= s40_val_n14;
    end
    always @(posedge \clk ) begin
        s41_val_n15 <= s40_val_n15;
    end
    always @(posedge \clk ) begin
        s41_val_n16 <= s40_val_n16;
    end
    always @(posedge \clk ) begin
        s41_val_n17 <= s40_val_n17;
    end
    always @(posedge \clk ) begin
        s41_val_n18 <= s40_val_n18;
    end
    always @(posedge \clk ) begin
        s41_val_n19 <= val_n19;
    end
    always @(posedge \clk ) begin
        \s42_val  <= \s41_val ;
    end
    always @(posedge \clk ) begin
        s42_val_n1 <= s41_val_n1;
    end
    always @(posedge \clk ) begin
        s42_val_n2 <= s41_val_n2;
    end
    always @(posedge \clk ) begin
        s42_val_n3 <= s41_val_n3;
    end
    always @(posedge \clk ) begin
        s42_val_n4 <= s41_val_n4;
    end
    always @(posedge \clk ) begin
        s42_val_n5 <= s41_val_n5;
    end
    always @(posedge \clk ) begin
        s42_val_n6 <= s41_val_n6;
    end
    always @(posedge \clk ) begin
        s42_val_n7 <= s41_val_n7;
    end
    always @(posedge \clk ) begin
        s42_val_n8 <= s41_val_n8;
    end
    always @(posedge \clk ) begin
        s42_val_n9 <= s41_val_n9;
    end
    always @(posedge \clk ) begin
        s42_val_n10 <= s41_val_n10;
    end
    always @(posedge \clk ) begin
        s42_val_n11 <= s41_val_n11;
    end
    always @(posedge \clk ) begin
        s42_val_n12 <= s41_val_n12;
    end
    always @(posedge \clk ) begin
        s42_val_n13 <= s41_val_n13;
    end
    always @(posedge \clk ) begin
        s42_val_n14 <= s41_val_n14;
    end
    always @(posedge \clk ) begin
        s42_val_n15 <= s41_val_n15;
    end
    always @(posedge \clk ) begin
        s42_val_n16 <= s41_val_n16;
    end
    always @(posedge \clk ) begin
        s42_val_n17 <= s41_val_n17;
    end
    always @(posedge \clk ) begin
        s42_val_n18 <= s41_val_n18;
    end
    always @(posedge \clk ) begin
        s42_val_n19 <= s41_val_n19;
    end
    always @(posedge \clk ) begin
        \s43_val  <= \s42_val ;
    end
    always @(posedge \clk ) begin
        s43_val_n1 <= s42_val_n1;
    end
    always @(posedge \clk ) begin
        s43_val_n2 <= s42_val_n2;
    end
    always @(posedge \clk ) begin
        s43_val_n3 <= s42_val_n3;
    end
    always @(posedge \clk ) begin
        s43_val_n4 <= s42_val_n4;
    end
    always @(posedge \clk ) begin
        s43_val_n5 <= s42_val_n5;
    end
    always @(posedge \clk ) begin
        s43_val_n6 <= s42_val_n6;
    end
    always @(posedge \clk ) begin
        s43_val_n7 <= s42_val_n7;
    end
    always @(posedge \clk ) begin
        s43_val_n8 <= s42_val_n8;
    end
    always @(posedge \clk ) begin
        s43_val_n9 <= s42_val_n9;
    end
    always @(posedge \clk ) begin
        s43_val_n10 <= s42_val_n10;
    end
    always @(posedge \clk ) begin
        s43_val_n11 <= s42_val_n11;
    end
    always @(posedge \clk ) begin
        s43_val_n12 <= s42_val_n12;
    end
    always @(posedge \clk ) begin
        s43_val_n13 <= s42_val_n13;
    end
    always @(posedge \clk ) begin
        s43_val_n14 <= s42_val_n14;
    end
    always @(posedge \clk ) begin
        s43_val_n15 <= s42_val_n15;
    end
    always @(posedge \clk ) begin
        s43_val_n16 <= s42_val_n16;
    end
    always @(posedge \clk ) begin
        s43_val_n17 <= s42_val_n17;
    end
    always @(posedge \clk ) begin
        s43_val_n18 <= s42_val_n18;
    end
    always @(posedge \clk ) begin
        s43_val_n19 <= s42_val_n19;
    end
    always @(posedge \clk ) begin
        s43_val_n20 <= val_n20;
    end
    always @(posedge \clk ) begin
        \s44_val  <= \s43_val ;
    end
    always @(posedge \clk ) begin
        s44_val_n1 <= s43_val_n1;
    end
    always @(posedge \clk ) begin
        s44_val_n2 <= s43_val_n2;
    end
    always @(posedge \clk ) begin
        s44_val_n3 <= s43_val_n3;
    end
    always @(posedge \clk ) begin
        s44_val_n4 <= s43_val_n4;
    end
    always @(posedge \clk ) begin
        s44_val_n5 <= s43_val_n5;
    end
    always @(posedge \clk ) begin
        s44_val_n6 <= s43_val_n6;
    end
    always @(posedge \clk ) begin
        s44_val_n7 <= s43_val_n7;
    end
    always @(posedge \clk ) begin
        s44_val_n8 <= s43_val_n8;
    end
    always @(posedge \clk ) begin
        s44_val_n9 <= s43_val_n9;
    end
    always @(posedge \clk ) begin
        s44_val_n10 <= s43_val_n10;
    end
    always @(posedge \clk ) begin
        s44_val_n11 <= s43_val_n11;
    end
    always @(posedge \clk ) begin
        s44_val_n12 <= s43_val_n12;
    end
    always @(posedge \clk ) begin
        s44_val_n13 <= s43_val_n13;
    end
    always @(posedge \clk ) begin
        s44_val_n14 <= s43_val_n14;
    end
    always @(posedge \clk ) begin
        s44_val_n15 <= s43_val_n15;
    end
    always @(posedge \clk ) begin
        s44_val_n16 <= s43_val_n16;
    end
    always @(posedge \clk ) begin
        s44_val_n17 <= s43_val_n17;
    end
    always @(posedge \clk ) begin
        s44_val_n18 <= s43_val_n18;
    end
    always @(posedge \clk ) begin
        s44_val_n19 <= s43_val_n19;
    end
    always @(posedge \clk ) begin
        s44_val_n20 <= s43_val_n20;
    end
    always @(posedge \clk ) begin
        \s45_val  <= \s44_val ;
    end
    always @(posedge \clk ) begin
        s45_val_n1 <= s44_val_n1;
    end
    always @(posedge \clk ) begin
        s45_val_n2 <= s44_val_n2;
    end
    always @(posedge \clk ) begin
        s45_val_n3 <= s44_val_n3;
    end
    always @(posedge \clk ) begin
        s45_val_n4 <= s44_val_n4;
    end
    always @(posedge \clk ) begin
        s45_val_n5 <= s44_val_n5;
    end
    always @(posedge \clk ) begin
        s45_val_n6 <= s44_val_n6;
    end
    always @(posedge \clk ) begin
        s45_val_n7 <= s44_val_n7;
    end
    always @(posedge \clk ) begin
        s45_val_n8 <= s44_val_n8;
    end
    always @(posedge \clk ) begin
        s45_val_n9 <= s44_val_n9;
    end
    always @(posedge \clk ) begin
        s45_val_n10 <= s44_val_n10;
    end
    always @(posedge \clk ) begin
        s45_val_n11 <= s44_val_n11;
    end
    always @(posedge \clk ) begin
        s45_val_n12 <= s44_val_n12;
    end
    always @(posedge \clk ) begin
        s45_val_n13 <= s44_val_n13;
    end
    always @(posedge \clk ) begin
        s45_val_n14 <= s44_val_n14;
    end
    always @(posedge \clk ) begin
        s45_val_n15 <= s44_val_n15;
    end
    always @(posedge \clk ) begin
        s45_val_n16 <= s44_val_n16;
    end
    always @(posedge \clk ) begin
        s45_val_n17 <= s44_val_n17;
    end
    always @(posedge \clk ) begin
        s45_val_n18 <= s44_val_n18;
    end
    always @(posedge \clk ) begin
        s45_val_n19 <= s44_val_n19;
    end
    always @(posedge \clk ) begin
        s45_val_n20 <= s44_val_n20;
    end
    always @(posedge \clk ) begin
        s45_val_n21 <= val_n21;
    end
    always @(posedge \clk ) begin
        \s46_val  <= \s45_val ;
    end
    always @(posedge \clk ) begin
        s46_val_n1 <= s45_val_n1;
    end
    always @(posedge \clk ) begin
        s46_val_n2 <= s45_val_n2;
    end
    always @(posedge \clk ) begin
        s46_val_n3 <= s45_val_n3;
    end
    always @(posedge \clk ) begin
        s46_val_n4 <= s45_val_n4;
    end
    always @(posedge \clk ) begin
        s46_val_n5 <= s45_val_n5;
    end
    always @(posedge \clk ) begin
        s46_val_n6 <= s45_val_n6;
    end
    always @(posedge \clk ) begin
        s46_val_n7 <= s45_val_n7;
    end
    always @(posedge \clk ) begin
        s46_val_n8 <= s45_val_n8;
    end
    always @(posedge \clk ) begin
        s46_val_n9 <= s45_val_n9;
    end
    always @(posedge \clk ) begin
        s46_val_n10 <= s45_val_n10;
    end
    always @(posedge \clk ) begin
        s46_val_n11 <= s45_val_n11;
    end
    always @(posedge \clk ) begin
        s46_val_n12 <= s45_val_n12;
    end
    always @(posedge \clk ) begin
        s46_val_n13 <= s45_val_n13;
    end
    always @(posedge \clk ) begin
        s46_val_n14 <= s45_val_n14;
    end
    always @(posedge \clk ) begin
        s46_val_n15 <= s45_val_n15;
    end
    always @(posedge \clk ) begin
        s46_val_n16 <= s45_val_n16;
    end
    always @(posedge \clk ) begin
        s46_val_n17 <= s45_val_n17;
    end
    always @(posedge \clk ) begin
        s46_val_n18 <= s45_val_n18;
    end
    always @(posedge \clk ) begin
        s46_val_n19 <= s45_val_n19;
    end
    always @(posedge \clk ) begin
        s46_val_n20 <= s45_val_n20;
    end
    always @(posedge \clk ) begin
        s46_val_n21 <= s45_val_n21;
    end
    always @(posedge \clk ) begin
        \s47_val  <= \s46_val ;
    end
    always @(posedge \clk ) begin
        s47_val_n1 <= s46_val_n1;
    end
    always @(posedge \clk ) begin
        s47_val_n2 <= s46_val_n2;
    end
    always @(posedge \clk ) begin
        s47_val_n3 <= s46_val_n3;
    end
    always @(posedge \clk ) begin
        s47_val_n4 <= s46_val_n4;
    end
    always @(posedge \clk ) begin
        s47_val_n5 <= s46_val_n5;
    end
    always @(posedge \clk ) begin
        s47_val_n6 <= s46_val_n6;
    end
    always @(posedge \clk ) begin
        s47_val_n7 <= s46_val_n7;
    end
    always @(posedge \clk ) begin
        s47_val_n8 <= s46_val_n8;
    end
    always @(posedge \clk ) begin
        s47_val_n9 <= s46_val_n9;
    end
    always @(posedge \clk ) begin
        s47_val_n10 <= s46_val_n10;
    end
    always @(posedge \clk ) begin
        s47_val_n11 <= s46_val_n11;
    end
    always @(posedge \clk ) begin
        s47_val_n12 <= s46_val_n12;
    end
    always @(posedge \clk ) begin
        s47_val_n13 <= s46_val_n13;
    end
    always @(posedge \clk ) begin
        s47_val_n14 <= s46_val_n14;
    end
    always @(posedge \clk ) begin
        s47_val_n15 <= s46_val_n15;
    end
    always @(posedge \clk ) begin
        s47_val_n16 <= s46_val_n16;
    end
    always @(posedge \clk ) begin
        s47_val_n17 <= s46_val_n17;
    end
    always @(posedge \clk ) begin
        s47_val_n18 <= s46_val_n18;
    end
    always @(posedge \clk ) begin
        s47_val_n19 <= s46_val_n19;
    end
    always @(posedge \clk ) begin
        s47_val_n20 <= s46_val_n20;
    end
    always @(posedge \clk ) begin
        s47_val_n21 <= s46_val_n21;
    end
    always @(posedge \clk ) begin
        s47_val_n22 <= val_n22;
    end
    always @(posedge \clk ) begin
        \s48_val  <= \s47_val ;
    end
    always @(posedge \clk ) begin
        s48_val_n1 <= s47_val_n1;
    end
    always @(posedge \clk ) begin
        s48_val_n2 <= s47_val_n2;
    end
    always @(posedge \clk ) begin
        s48_val_n3 <= s47_val_n3;
    end
    always @(posedge \clk ) begin
        s48_val_n4 <= s47_val_n4;
    end
    always @(posedge \clk ) begin
        s48_val_n5 <= s47_val_n5;
    end
    always @(posedge \clk ) begin
        s48_val_n6 <= s47_val_n6;
    end
    always @(posedge \clk ) begin
        s48_val_n7 <= s47_val_n7;
    end
    always @(posedge \clk ) begin
        s48_val_n8 <= s47_val_n8;
    end
    always @(posedge \clk ) begin
        s48_val_n9 <= s47_val_n9;
    end
    always @(posedge \clk ) begin
        s48_val_n10 <= s47_val_n10;
    end
    always @(posedge \clk ) begin
        s48_val_n11 <= s47_val_n11;
    end
    always @(posedge \clk ) begin
        s48_val_n12 <= s47_val_n12;
    end
    always @(posedge \clk ) begin
        s48_val_n13 <= s47_val_n13;
    end
    always @(posedge \clk ) begin
        s48_val_n14 <= s47_val_n14;
    end
    always @(posedge \clk ) begin
        s48_val_n15 <= s47_val_n15;
    end
    always @(posedge \clk ) begin
        s48_val_n16 <= s47_val_n16;
    end
    always @(posedge \clk ) begin
        s48_val_n17 <= s47_val_n17;
    end
    always @(posedge \clk ) begin
        s48_val_n18 <= s47_val_n18;
    end
    always @(posedge \clk ) begin
        s48_val_n19 <= s47_val_n19;
    end
    always @(posedge \clk ) begin
        s48_val_n20 <= s47_val_n20;
    end
    always @(posedge \clk ) begin
        s48_val_n21 <= s47_val_n21;
    end
    always @(posedge \clk ) begin
        s48_val_n22 <= s47_val_n22;
    end
    always @(posedge \clk ) begin
        \s49_val  <= \s48_val ;
    end
    always @(posedge \clk ) begin
        s49_val_n1 <= s48_val_n1;
    end
    always @(posedge \clk ) begin
        s49_val_n2 <= s48_val_n2;
    end
    always @(posedge \clk ) begin
        s49_val_n3 <= s48_val_n3;
    end
    always @(posedge \clk ) begin
        s49_val_n4 <= s48_val_n4;
    end
    always @(posedge \clk ) begin
        s49_val_n5 <= s48_val_n5;
    end
    always @(posedge \clk ) begin
        s49_val_n6 <= s48_val_n6;
    end
    always @(posedge \clk ) begin
        s49_val_n7 <= s48_val_n7;
    end
    always @(posedge \clk ) begin
        s49_val_n8 <= s48_val_n8;
    end
    always @(posedge \clk ) begin
        s49_val_n9 <= s48_val_n9;
    end
    always @(posedge \clk ) begin
        s49_val_n10 <= s48_val_n10;
    end
    always @(posedge \clk ) begin
        s49_val_n11 <= s48_val_n11;
    end
    always @(posedge \clk ) begin
        s49_val_n12 <= s48_val_n12;
    end
    always @(posedge \clk ) begin
        s49_val_n13 <= s48_val_n13;
    end
    always @(posedge \clk ) begin
        s49_val_n14 <= s48_val_n14;
    end
    always @(posedge \clk ) begin
        s49_val_n15 <= s48_val_n15;
    end
    always @(posedge \clk ) begin
        s49_val_n16 <= s48_val_n16;
    end
    always @(posedge \clk ) begin
        s49_val_n17 <= s48_val_n17;
    end
    always @(posedge \clk ) begin
        s49_val_n18 <= s48_val_n18;
    end
    always @(posedge \clk ) begin
        s49_val_n19 <= s48_val_n19;
    end
    always @(posedge \clk ) begin
        s49_val_n20 <= s48_val_n20;
    end
    always @(posedge \clk ) begin
        s49_val_n21 <= s48_val_n21;
    end
    always @(posedge \clk ) begin
        s49_val_n22 <= s48_val_n22;
    end
    always @(posedge \clk ) begin
        s49_val_n23 <= val_n23;
    end
    always @(posedge \clk ) begin
        \s50_val  <= \s49_val ;
    end
    always @(posedge \clk ) begin
        s50_val_n1 <= s49_val_n1;
    end
    always @(posedge \clk ) begin
        s50_val_n2 <= s49_val_n2;
    end
    always @(posedge \clk ) begin
        s50_val_n3 <= s49_val_n3;
    end
    always @(posedge \clk ) begin
        s50_val_n4 <= s49_val_n4;
    end
    always @(posedge \clk ) begin
        s50_val_n5 <= s49_val_n5;
    end
    always @(posedge \clk ) begin
        s50_val_n6 <= s49_val_n6;
    end
    always @(posedge \clk ) begin
        s50_val_n7 <= s49_val_n7;
    end
    always @(posedge \clk ) begin
        s50_val_n8 <= s49_val_n8;
    end
    always @(posedge \clk ) begin
        s50_val_n9 <= s49_val_n9;
    end
    always @(posedge \clk ) begin
        s50_val_n10 <= s49_val_n10;
    end
    always @(posedge \clk ) begin
        s50_val_n11 <= s49_val_n11;
    end
    always @(posedge \clk ) begin
        s50_val_n12 <= s49_val_n12;
    end
    always @(posedge \clk ) begin
        s50_val_n13 <= s49_val_n13;
    end
    always @(posedge \clk ) begin
        s50_val_n14 <= s49_val_n14;
    end
    always @(posedge \clk ) begin
        s50_val_n15 <= s49_val_n15;
    end
    always @(posedge \clk ) begin
        s50_val_n16 <= s49_val_n16;
    end
    always @(posedge \clk ) begin
        s50_val_n17 <= s49_val_n17;
    end
    always @(posedge \clk ) begin
        s50_val_n18 <= s49_val_n18;
    end
    always @(posedge \clk ) begin
        s50_val_n19 <= s49_val_n19;
    end
    always @(posedge \clk ) begin
        s50_val_n20 <= s49_val_n20;
    end
    always @(posedge \clk ) begin
        s50_val_n21 <= s49_val_n21;
    end
    always @(posedge \clk ) begin
        s50_val_n22 <= s49_val_n22;
    end
    always @(posedge \clk ) begin
        s50_val_n23 <= s49_val_n23;
    end
    always @(posedge \clk ) begin
        \s51_val  <= \s50_val ;
    end
    always @(posedge \clk ) begin
        s51_val_n1 <= s50_val_n1;
    end
    always @(posedge \clk ) begin
        s51_val_n2 <= s50_val_n2;
    end
    always @(posedge \clk ) begin
        s51_val_n3 <= s50_val_n3;
    end
    always @(posedge \clk ) begin
        s51_val_n4 <= s50_val_n4;
    end
    always @(posedge \clk ) begin
        s51_val_n5 <= s50_val_n5;
    end
    always @(posedge \clk ) begin
        s51_val_n6 <= s50_val_n6;
    end
    always @(posedge \clk ) begin
        s51_val_n7 <= s50_val_n7;
    end
    always @(posedge \clk ) begin
        s51_val_n8 <= s50_val_n8;
    end
    always @(posedge \clk ) begin
        s51_val_n9 <= s50_val_n9;
    end
    always @(posedge \clk ) begin
        s51_val_n10 <= s50_val_n10;
    end
    always @(posedge \clk ) begin
        s51_val_n11 <= s50_val_n11;
    end
    always @(posedge \clk ) begin
        s51_val_n12 <= s50_val_n12;
    end
    always @(posedge \clk ) begin
        s51_val_n13 <= s50_val_n13;
    end
    always @(posedge \clk ) begin
        s51_val_n14 <= s50_val_n14;
    end
    always @(posedge \clk ) begin
        s51_val_n15 <= s50_val_n15;
    end
    always @(posedge \clk ) begin
        s51_val_n16 <= s50_val_n16;
    end
    always @(posedge \clk ) begin
        s51_val_n17 <= s50_val_n17;
    end
    always @(posedge \clk ) begin
        s51_val_n18 <= s50_val_n18;
    end
    always @(posedge \clk ) begin
        s51_val_n19 <= s50_val_n19;
    end
    always @(posedge \clk ) begin
        s51_val_n20 <= s50_val_n20;
    end
    always @(posedge \clk ) begin
        s51_val_n21 <= s50_val_n21;
    end
    always @(posedge \clk ) begin
        s51_val_n22 <= s50_val_n22;
    end
    always @(posedge \clk ) begin
        s51_val_n23 <= s50_val_n23;
    end
    always @(posedge \clk ) begin
        s51_val_n24 <= val_n24;
    end
    always @(posedge \clk ) begin
        \s52_val  <= \s51_val ;
    end
    always @(posedge \clk ) begin
        s52_val_n1 <= s51_val_n1;
    end
    always @(posedge \clk ) begin
        s52_val_n2 <= s51_val_n2;
    end
    always @(posedge \clk ) begin
        s52_val_n3 <= s51_val_n3;
    end
    always @(posedge \clk ) begin
        s52_val_n4 <= s51_val_n4;
    end
    always @(posedge \clk ) begin
        s52_val_n5 <= s51_val_n5;
    end
    always @(posedge \clk ) begin
        s52_val_n6 <= s51_val_n6;
    end
    always @(posedge \clk ) begin
        s52_val_n7 <= s51_val_n7;
    end
    always @(posedge \clk ) begin
        s52_val_n8 <= s51_val_n8;
    end
    always @(posedge \clk ) begin
        s52_val_n9 <= s51_val_n9;
    end
    always @(posedge \clk ) begin
        s52_val_n10 <= s51_val_n10;
    end
    always @(posedge \clk ) begin
        s52_val_n11 <= s51_val_n11;
    end
    always @(posedge \clk ) begin
        s52_val_n12 <= s51_val_n12;
    end
    always @(posedge \clk ) begin
        s52_val_n13 <= s51_val_n13;
    end
    always @(posedge \clk ) begin
        s52_val_n14 <= s51_val_n14;
    end
    always @(posedge \clk ) begin
        s52_val_n15 <= s51_val_n15;
    end
    always @(posedge \clk ) begin
        s52_val_n16 <= s51_val_n16;
    end
    always @(posedge \clk ) begin
        s52_val_n17 <= s51_val_n17;
    end
    always @(posedge \clk ) begin
        s52_val_n18 <= s51_val_n18;
    end
    always @(posedge \clk ) begin
        s52_val_n19 <= s51_val_n19;
    end
    always @(posedge \clk ) begin
        s52_val_n20 <= s51_val_n20;
    end
    always @(posedge \clk ) begin
        s52_val_n21 <= s51_val_n21;
    end
    always @(posedge \clk ) begin
        s52_val_n22 <= s51_val_n22;
    end
    always @(posedge \clk ) begin
        s52_val_n23 <= s51_val_n23;
    end
    always @(posedge \clk ) begin
        s52_val_n24 <= s51_val_n24;
    end
    always @(posedge \clk ) begin
        \s53_val  <= \s52_val ;
    end
    always @(posedge \clk ) begin
        s53_val_n1 <= s52_val_n1;
    end
    always @(posedge \clk ) begin
        s53_val_n2 <= s52_val_n2;
    end
    always @(posedge \clk ) begin
        s53_val_n3 <= s52_val_n3;
    end
    always @(posedge \clk ) begin
        s53_val_n4 <= s52_val_n4;
    end
    always @(posedge \clk ) begin
        s53_val_n5 <= s52_val_n5;
    end
    always @(posedge \clk ) begin
        s53_val_n6 <= s52_val_n6;
    end
    always @(posedge \clk ) begin
        s53_val_n7 <= s52_val_n7;
    end
    always @(posedge \clk ) begin
        s53_val_n8 <= s52_val_n8;
    end
    always @(posedge \clk ) begin
        s53_val_n9 <= s52_val_n9;
    end
    always @(posedge \clk ) begin
        s53_val_n10 <= s52_val_n10;
    end
    always @(posedge \clk ) begin
        s53_val_n11 <= s52_val_n11;
    end
    always @(posedge \clk ) begin
        s53_val_n12 <= s52_val_n12;
    end
    always @(posedge \clk ) begin
        s53_val_n13 <= s52_val_n13;
    end
    always @(posedge \clk ) begin
        s53_val_n14 <= s52_val_n14;
    end
    always @(posedge \clk ) begin
        s53_val_n15 <= s52_val_n15;
    end
    always @(posedge \clk ) begin
        s53_val_n16 <= s52_val_n16;
    end
    always @(posedge \clk ) begin
        s53_val_n17 <= s52_val_n17;
    end
    always @(posedge \clk ) begin
        s53_val_n18 <= s52_val_n18;
    end
    always @(posedge \clk ) begin
        s53_val_n19 <= s52_val_n19;
    end
    always @(posedge \clk ) begin
        s53_val_n20 <= s52_val_n20;
    end
    always @(posedge \clk ) begin
        s53_val_n21 <= s52_val_n21;
    end
    always @(posedge \clk ) begin
        s53_val_n22 <= s52_val_n22;
    end
    always @(posedge \clk ) begin
        s53_val_n23 <= s52_val_n23;
    end
    always @(posedge \clk ) begin
        s53_val_n24 <= s52_val_n24;
    end
    always @(posedge \clk ) begin
        s53_val_n25 <= val_n25;
    end
    always @(posedge \clk ) begin
        \s54_val  <= \s53_val ;
    end
    always @(posedge \clk ) begin
        s54_val_n1 <= s53_val_n1;
    end
    always @(posedge \clk ) begin
        s54_val_n2 <= s53_val_n2;
    end
    always @(posedge \clk ) begin
        s54_val_n3 <= s53_val_n3;
    end
    always @(posedge \clk ) begin
        s54_val_n4 <= s53_val_n4;
    end
    always @(posedge \clk ) begin
        s54_val_n5 <= s53_val_n5;
    end
    always @(posedge \clk ) begin
        s54_val_n6 <= s53_val_n6;
    end
    always @(posedge \clk ) begin
        s54_val_n7 <= s53_val_n7;
    end
    always @(posedge \clk ) begin
        s54_val_n8 <= s53_val_n8;
    end
    always @(posedge \clk ) begin
        s54_val_n9 <= s53_val_n9;
    end
    always @(posedge \clk ) begin
        s54_val_n10 <= s53_val_n10;
    end
    always @(posedge \clk ) begin
        s54_val_n11 <= s53_val_n11;
    end
    always @(posedge \clk ) begin
        s54_val_n12 <= s53_val_n12;
    end
    always @(posedge \clk ) begin
        s54_val_n13 <= s53_val_n13;
    end
    always @(posedge \clk ) begin
        s54_val_n14 <= s53_val_n14;
    end
    always @(posedge \clk ) begin
        s54_val_n15 <= s53_val_n15;
    end
    always @(posedge \clk ) begin
        s54_val_n16 <= s53_val_n16;
    end
    always @(posedge \clk ) begin
        s54_val_n17 <= s53_val_n17;
    end
    always @(posedge \clk ) begin
        s54_val_n18 <= s53_val_n18;
    end
    always @(posedge \clk ) begin
        s54_val_n19 <= s53_val_n19;
    end
    always @(posedge \clk ) begin
        s54_val_n20 <= s53_val_n20;
    end
    always @(posedge \clk ) begin
        s54_val_n21 <= s53_val_n21;
    end
    always @(posedge \clk ) begin
        s54_val_n22 <= s53_val_n22;
    end
    always @(posedge \clk ) begin
        s54_val_n23 <= s53_val_n23;
    end
    always @(posedge \clk ) begin
        s54_val_n24 <= s53_val_n24;
    end
    always @(posedge \clk ) begin
        s54_val_n25 <= s53_val_n25;
    end
    always @(posedge \clk ) begin
        \s55_val  <= \s54_val ;
    end
    always @(posedge \clk ) begin
        s55_val_n1 <= s54_val_n1;
    end
    always @(posedge \clk ) begin
        s55_val_n2 <= s54_val_n2;
    end
    always @(posedge \clk ) begin
        s55_val_n3 <= s54_val_n3;
    end
    always @(posedge \clk ) begin
        s55_val_n4 <= s54_val_n4;
    end
    always @(posedge \clk ) begin
        s55_val_n5 <= s54_val_n5;
    end
    always @(posedge \clk ) begin
        s55_val_n6 <= s54_val_n6;
    end
    always @(posedge \clk ) begin
        s55_val_n7 <= s54_val_n7;
    end
    always @(posedge \clk ) begin
        s55_val_n8 <= s54_val_n8;
    end
    always @(posedge \clk ) begin
        s55_val_n9 <= s54_val_n9;
    end
    always @(posedge \clk ) begin
        s55_val_n10 <= s54_val_n10;
    end
    always @(posedge \clk ) begin
        s55_val_n11 <= s54_val_n11;
    end
    always @(posedge \clk ) begin
        s55_val_n12 <= s54_val_n12;
    end
    always @(posedge \clk ) begin
        s55_val_n13 <= s54_val_n13;
    end
    always @(posedge \clk ) begin
        s55_val_n14 <= s54_val_n14;
    end
    always @(posedge \clk ) begin
        s55_val_n15 <= s54_val_n15;
    end
    always @(posedge \clk ) begin
        s55_val_n16 <= s54_val_n16;
    end
    always @(posedge \clk ) begin
        s55_val_n17 <= s54_val_n17;
    end
    always @(posedge \clk ) begin
        s55_val_n18 <= s54_val_n18;
    end
    always @(posedge \clk ) begin
        s55_val_n19 <= s54_val_n19;
    end
    always @(posedge \clk ) begin
        s55_val_n20 <= s54_val_n20;
    end
    always @(posedge \clk ) begin
        s55_val_n21 <= s54_val_n21;
    end
    always @(posedge \clk ) begin
        s55_val_n22 <= s54_val_n22;
    end
    always @(posedge \clk ) begin
        s55_val_n23 <= s54_val_n23;
    end
    always @(posedge \clk ) begin
        s55_val_n24 <= s54_val_n24;
    end
    always @(posedge \clk ) begin
        s55_val_n25 <= s54_val_n25;
    end
    always @(posedge \clk ) begin
        s55_val_n26 <= val_n26;
    end
    always @(posedge \clk ) begin
        \s56_val  <= \s55_val ;
    end
    always @(posedge \clk ) begin
        s56_val_n1 <= s55_val_n1;
    end
    always @(posedge \clk ) begin
        s56_val_n2 <= s55_val_n2;
    end
    always @(posedge \clk ) begin
        s56_val_n3 <= s55_val_n3;
    end
    always @(posedge \clk ) begin
        s56_val_n4 <= s55_val_n4;
    end
    always @(posedge \clk ) begin
        s56_val_n5 <= s55_val_n5;
    end
    always @(posedge \clk ) begin
        s56_val_n6 <= s55_val_n6;
    end
    always @(posedge \clk ) begin
        s56_val_n7 <= s55_val_n7;
    end
    always @(posedge \clk ) begin
        s56_val_n8 <= s55_val_n8;
    end
    always @(posedge \clk ) begin
        s56_val_n9 <= s55_val_n9;
    end
    always @(posedge \clk ) begin
        s56_val_n10 <= s55_val_n10;
    end
    always @(posedge \clk ) begin
        s56_val_n11 <= s55_val_n11;
    end
    always @(posedge \clk ) begin
        s56_val_n12 <= s55_val_n12;
    end
    always @(posedge \clk ) begin
        s56_val_n13 <= s55_val_n13;
    end
    always @(posedge \clk ) begin
        s56_val_n14 <= s55_val_n14;
    end
    always @(posedge \clk ) begin
        s56_val_n15 <= s55_val_n15;
    end
    always @(posedge \clk ) begin
        s56_val_n16 <= s55_val_n16;
    end
    always @(posedge \clk ) begin
        s56_val_n17 <= s55_val_n17;
    end
    always @(posedge \clk ) begin
        s56_val_n18 <= s55_val_n18;
    end
    always @(posedge \clk ) begin
        s56_val_n19 <= s55_val_n19;
    end
    always @(posedge \clk ) begin
        s56_val_n20 <= s55_val_n20;
    end
    always @(posedge \clk ) begin
        s56_val_n21 <= s55_val_n21;
    end
    always @(posedge \clk ) begin
        s56_val_n22 <= s55_val_n22;
    end
    always @(posedge \clk ) begin
        s56_val_n23 <= s55_val_n23;
    end
    always @(posedge \clk ) begin
        s56_val_n24 <= s55_val_n24;
    end
    always @(posedge \clk ) begin
        s56_val_n25 <= s55_val_n25;
    end
    always @(posedge \clk ) begin
        s56_val_n26 <= s55_val_n26;
    end
    always @(posedge \clk ) begin
        \s57_val  <= \s56_val ;
    end
    always @(posedge \clk ) begin
        s57_val_n1 <= s56_val_n1;
    end
    always @(posedge \clk ) begin
        s57_val_n2 <= s56_val_n2;
    end
    always @(posedge \clk ) begin
        s57_val_n3 <= s56_val_n3;
    end
    always @(posedge \clk ) begin
        s57_val_n4 <= s56_val_n4;
    end
    always @(posedge \clk ) begin
        s57_val_n5 <= s56_val_n5;
    end
    always @(posedge \clk ) begin
        s57_val_n6 <= s56_val_n6;
    end
    always @(posedge \clk ) begin
        s57_val_n7 <= s56_val_n7;
    end
    always @(posedge \clk ) begin
        s57_val_n8 <= s56_val_n8;
    end
    always @(posedge \clk ) begin
        s57_val_n9 <= s56_val_n9;
    end
    always @(posedge \clk ) begin
        s57_val_n10 <= s56_val_n10;
    end
    always @(posedge \clk ) begin
        s57_val_n11 <= s56_val_n11;
    end
    always @(posedge \clk ) begin
        s57_val_n12 <= s56_val_n12;
    end
    always @(posedge \clk ) begin
        s57_val_n13 <= s56_val_n13;
    end
    always @(posedge \clk ) begin
        s57_val_n14 <= s56_val_n14;
    end
    always @(posedge \clk ) begin
        s57_val_n15 <= s56_val_n15;
    end
    always @(posedge \clk ) begin
        s57_val_n16 <= s56_val_n16;
    end
    always @(posedge \clk ) begin
        s57_val_n17 <= s56_val_n17;
    end
    always @(posedge \clk ) begin
        s57_val_n18 <= s56_val_n18;
    end
    always @(posedge \clk ) begin
        s57_val_n19 <= s56_val_n19;
    end
    always @(posedge \clk ) begin
        s57_val_n20 <= s56_val_n20;
    end
    always @(posedge \clk ) begin
        s57_val_n21 <= s56_val_n21;
    end
    always @(posedge \clk ) begin
        s57_val_n22 <= s56_val_n22;
    end
    always @(posedge \clk ) begin
        s57_val_n23 <= s56_val_n23;
    end
    always @(posedge \clk ) begin
        s57_val_n24 <= s56_val_n24;
    end
    always @(posedge \clk ) begin
        s57_val_n25 <= s56_val_n25;
    end
    always @(posedge \clk ) begin
        s57_val_n26 <= s56_val_n26;
    end
    always @(posedge \clk ) begin
        s57_val_n27 <= val_n27;
    end
    always @(posedge \clk ) begin
        \s58_val  <= \s57_val ;
    end
    always @(posedge \clk ) begin
        s58_val_n1 <= s57_val_n1;
    end
    always @(posedge \clk ) begin
        s58_val_n2 <= s57_val_n2;
    end
    always @(posedge \clk ) begin
        s58_val_n3 <= s57_val_n3;
    end
    always @(posedge \clk ) begin
        s58_val_n4 <= s57_val_n4;
    end
    always @(posedge \clk ) begin
        s58_val_n5 <= s57_val_n5;
    end
    always @(posedge \clk ) begin
        s58_val_n6 <= s57_val_n6;
    end
    always @(posedge \clk ) begin
        s58_val_n7 <= s57_val_n7;
    end
    always @(posedge \clk ) begin
        s58_val_n8 <= s57_val_n8;
    end
    always @(posedge \clk ) begin
        s58_val_n9 <= s57_val_n9;
    end
    always @(posedge \clk ) begin
        s58_val_n10 <= s57_val_n10;
    end
    always @(posedge \clk ) begin
        s58_val_n11 <= s57_val_n11;
    end
    always @(posedge \clk ) begin
        s58_val_n12 <= s57_val_n12;
    end
    always @(posedge \clk ) begin
        s58_val_n13 <= s57_val_n13;
    end
    always @(posedge \clk ) begin
        s58_val_n14 <= s57_val_n14;
    end
    always @(posedge \clk ) begin
        s58_val_n15 <= s57_val_n15;
    end
    always @(posedge \clk ) begin
        s58_val_n16 <= s57_val_n16;
    end
    always @(posedge \clk ) begin
        s58_val_n17 <= s57_val_n17;
    end
    always @(posedge \clk ) begin
        s58_val_n18 <= s57_val_n18;
    end
    always @(posedge \clk ) begin
        s58_val_n19 <= s57_val_n19;
    end
    always @(posedge \clk ) begin
        s58_val_n20 <= s57_val_n20;
    end
    always @(posedge \clk ) begin
        s58_val_n21 <= s57_val_n21;
    end
    always @(posedge \clk ) begin
        s58_val_n22 <= s57_val_n22;
    end
    always @(posedge \clk ) begin
        s58_val_n23 <= s57_val_n23;
    end
    always @(posedge \clk ) begin
        s58_val_n24 <= s57_val_n24;
    end
    always @(posedge \clk ) begin
        s58_val_n25 <= s57_val_n25;
    end
    always @(posedge \clk ) begin
        s58_val_n26 <= s57_val_n26;
    end
    always @(posedge \clk ) begin
        s58_val_n27 <= s57_val_n27;
    end
    always @(posedge \clk ) begin
        \s59_val  <= \s58_val ;
    end
    always @(posedge \clk ) begin
        s59_val_n1 <= s58_val_n1;
    end
    always @(posedge \clk ) begin
        s59_val_n2 <= s58_val_n2;
    end
    always @(posedge \clk ) begin
        s59_val_n3 <= s58_val_n3;
    end
    always @(posedge \clk ) begin
        s59_val_n4 <= s58_val_n4;
    end
    always @(posedge \clk ) begin
        s59_val_n5 <= s58_val_n5;
    end
    always @(posedge \clk ) begin
        s59_val_n6 <= s58_val_n6;
    end
    always @(posedge \clk ) begin
        s59_val_n7 <= s58_val_n7;
    end
    always @(posedge \clk ) begin
        s59_val_n8 <= s58_val_n8;
    end
    always @(posedge \clk ) begin
        s59_val_n9 <= s58_val_n9;
    end
    always @(posedge \clk ) begin
        s59_val_n10 <= s58_val_n10;
    end
    always @(posedge \clk ) begin
        s59_val_n11 <= s58_val_n11;
    end
    always @(posedge \clk ) begin
        s59_val_n12 <= s58_val_n12;
    end
    always @(posedge \clk ) begin
        s59_val_n13 <= s58_val_n13;
    end
    always @(posedge \clk ) begin
        s59_val_n14 <= s58_val_n14;
    end
    always @(posedge \clk ) begin
        s59_val_n15 <= s58_val_n15;
    end
    always @(posedge \clk ) begin
        s59_val_n16 <= s58_val_n16;
    end
    always @(posedge \clk ) begin
        s59_val_n17 <= s58_val_n17;
    end
    always @(posedge \clk ) begin
        s59_val_n18 <= s58_val_n18;
    end
    always @(posedge \clk ) begin
        s59_val_n19 <= s58_val_n19;
    end
    always @(posedge \clk ) begin
        s59_val_n20 <= s58_val_n20;
    end
    always @(posedge \clk ) begin
        s59_val_n21 <= s58_val_n21;
    end
    always @(posedge \clk ) begin
        s59_val_n22 <= s58_val_n22;
    end
    always @(posedge \clk ) begin
        s59_val_n23 <= s58_val_n23;
    end
    always @(posedge \clk ) begin
        s59_val_n24 <= s58_val_n24;
    end
    always @(posedge \clk ) begin
        s59_val_n25 <= s58_val_n25;
    end
    always @(posedge \clk ) begin
        s59_val_n26 <= s58_val_n26;
    end
    always @(posedge \clk ) begin
        s59_val_n27 <= s58_val_n27;
    end
    always @(posedge \clk ) begin
        s59_val_n28 <= val_n28;
    end
    always @(posedge \clk ) begin
        \s60_val  <= \s59_val ;
    end
    always @(posedge \clk ) begin
        s60_val_n1 <= s59_val_n1;
    end
    always @(posedge \clk ) begin
        s60_val_n2 <= s59_val_n2;
    end
    always @(posedge \clk ) begin
        s60_val_n3 <= s59_val_n3;
    end
    always @(posedge \clk ) begin
        s60_val_n4 <= s59_val_n4;
    end
    always @(posedge \clk ) begin
        s60_val_n5 <= s59_val_n5;
    end
    always @(posedge \clk ) begin
        s60_val_n6 <= s59_val_n6;
    end
    always @(posedge \clk ) begin
        s60_val_n7 <= s59_val_n7;
    end
    always @(posedge \clk ) begin
        s60_val_n8 <= s59_val_n8;
    end
    always @(posedge \clk ) begin
        s60_val_n9 <= s59_val_n9;
    end
    always @(posedge \clk ) begin
        s60_val_n10 <= s59_val_n10;
    end
    always @(posedge \clk ) begin
        s60_val_n11 <= s59_val_n11;
    end
    always @(posedge \clk ) begin
        s60_val_n12 <= s59_val_n12;
    end
    always @(posedge \clk ) begin
        s60_val_n13 <= s59_val_n13;
    end
    always @(posedge \clk ) begin
        s60_val_n14 <= s59_val_n14;
    end
    always @(posedge \clk ) begin
        s60_val_n15 <= s59_val_n15;
    end
    always @(posedge \clk ) begin
        s60_val_n16 <= s59_val_n16;
    end
    always @(posedge \clk ) begin
        s60_val_n17 <= s59_val_n17;
    end
    always @(posedge \clk ) begin
        s60_val_n18 <= s59_val_n18;
    end
    always @(posedge \clk ) begin
        s60_val_n19 <= s59_val_n19;
    end
    always @(posedge \clk ) begin
        s60_val_n20 <= s59_val_n20;
    end
    always @(posedge \clk ) begin
        s60_val_n21 <= s59_val_n21;
    end
    always @(posedge \clk ) begin
        s60_val_n22 <= s59_val_n22;
    end
    always @(posedge \clk ) begin
        s60_val_n23 <= s59_val_n23;
    end
    always @(posedge \clk ) begin
        s60_val_n24 <= s59_val_n24;
    end
    always @(posedge \clk ) begin
        s60_val_n25 <= s59_val_n25;
    end
    always @(posedge \clk ) begin
        s60_val_n26 <= s59_val_n26;
    end
    always @(posedge \clk ) begin
        s60_val_n27 <= s59_val_n27;
    end
    always @(posedge \clk ) begin
        s60_val_n28 <= s59_val_n28;
    end
    always @(posedge \clk ) begin
        \s61_val  <= \s60_val ;
    end
    always @(posedge \clk ) begin
        s61_val_n1 <= s60_val_n1;
    end
    always @(posedge \clk ) begin
        s61_val_n2 <= s60_val_n2;
    end
    always @(posedge \clk ) begin
        s61_val_n3 <= s60_val_n3;
    end
    always @(posedge \clk ) begin
        s61_val_n4 <= s60_val_n4;
    end
    always @(posedge \clk ) begin
        s61_val_n5 <= s60_val_n5;
    end
    always @(posedge \clk ) begin
        s61_val_n6 <= s60_val_n6;
    end
    always @(posedge \clk ) begin
        s61_val_n7 <= s60_val_n7;
    end
    always @(posedge \clk ) begin
        s61_val_n8 <= s60_val_n8;
    end
    always @(posedge \clk ) begin
        s61_val_n9 <= s60_val_n9;
    end
    always @(posedge \clk ) begin
        s61_val_n10 <= s60_val_n10;
    end
    always @(posedge \clk ) begin
        s61_val_n11 <= s60_val_n11;
    end
    always @(posedge \clk ) begin
        s61_val_n12 <= s60_val_n12;
    end
    always @(posedge \clk ) begin
        s61_val_n13 <= s60_val_n13;
    end
    always @(posedge \clk ) begin
        s61_val_n14 <= s60_val_n14;
    end
    always @(posedge \clk ) begin
        s61_val_n15 <= s60_val_n15;
    end
    always @(posedge \clk ) begin
        s61_val_n16 <= s60_val_n16;
    end
    always @(posedge \clk ) begin
        s61_val_n17 <= s60_val_n17;
    end
    always @(posedge \clk ) begin
        s61_val_n18 <= s60_val_n18;
    end
    always @(posedge \clk ) begin
        s61_val_n19 <= s60_val_n19;
    end
    always @(posedge \clk ) begin
        s61_val_n20 <= s60_val_n20;
    end
    always @(posedge \clk ) begin
        s61_val_n21 <= s60_val_n21;
    end
    always @(posedge \clk ) begin
        s61_val_n22 <= s60_val_n22;
    end
    always @(posedge \clk ) begin
        s61_val_n23 <= s60_val_n23;
    end
    always @(posedge \clk ) begin
        s61_val_n24 <= s60_val_n24;
    end
    always @(posedge \clk ) begin
        s61_val_n25 <= s60_val_n25;
    end
    always @(posedge \clk ) begin
        s61_val_n26 <= s60_val_n26;
    end
    always @(posedge \clk ) begin
        s61_val_n27 <= s60_val_n27;
    end
    always @(posedge \clk ) begin
        s61_val_n28 <= s60_val_n28;
    end
    always @(posedge \clk ) begin
        s61_val_n29 <= val_n29;
    end
    always @(posedge \clk ) begin
        \s62_val  <= \s61_val ;
    end
    always @(posedge \clk ) begin
        s62_val_n1 <= s61_val_n1;
    end
    always @(posedge \clk ) begin
        s62_val_n2 <= s61_val_n2;
    end
    always @(posedge \clk ) begin
        s62_val_n3 <= s61_val_n3;
    end
    always @(posedge \clk ) begin
        s62_val_n4 <= s61_val_n4;
    end
    always @(posedge \clk ) begin
        s62_val_n5 <= s61_val_n5;
    end
    always @(posedge \clk ) begin
        s62_val_n6 <= s61_val_n6;
    end
    always @(posedge \clk ) begin
        s62_val_n7 <= s61_val_n7;
    end
    always @(posedge \clk ) begin
        s62_val_n8 <= s61_val_n8;
    end
    always @(posedge \clk ) begin
        s62_val_n9 <= s61_val_n9;
    end
    always @(posedge \clk ) begin
        s62_val_n10 <= s61_val_n10;
    end
    always @(posedge \clk ) begin
        s62_val_n11 <= s61_val_n11;
    end
    always @(posedge \clk ) begin
        s62_val_n12 <= s61_val_n12;
    end
    always @(posedge \clk ) begin
        s62_val_n13 <= s61_val_n13;
    end
    always @(posedge \clk ) begin
        s62_val_n14 <= s61_val_n14;
    end
    always @(posedge \clk ) begin
        s62_val_n15 <= s61_val_n15;
    end
    always @(posedge \clk ) begin
        s62_val_n16 <= s61_val_n16;
    end
    always @(posedge \clk ) begin
        s62_val_n17 <= s61_val_n17;
    end
    always @(posedge \clk ) begin
        s62_val_n18 <= s61_val_n18;
    end
    always @(posedge \clk ) begin
        s62_val_n19 <= s61_val_n19;
    end
    always @(posedge \clk ) begin
        s62_val_n20 <= s61_val_n20;
    end
    always @(posedge \clk ) begin
        s62_val_n21 <= s61_val_n21;
    end
    always @(posedge \clk ) begin
        s62_val_n22 <= s61_val_n22;
    end
    always @(posedge \clk ) begin
        s62_val_n23 <= s61_val_n23;
    end
    always @(posedge \clk ) begin
        s62_val_n24 <= s61_val_n24;
    end
    always @(posedge \clk ) begin
        s62_val_n25 <= s61_val_n25;
    end
    always @(posedge \clk ) begin
        s62_val_n26 <= s61_val_n26;
    end
    always @(posedge \clk ) begin
        s62_val_n27 <= s61_val_n27;
    end
    always @(posedge \clk ) begin
        s62_val_n28 <= s61_val_n28;
    end
    always @(posedge \clk ) begin
        s62_val_n29 <= s61_val_n29;
    end
    always @(posedge \clk ) begin
        \s63_val  <= \s62_val ;
    end
    always @(posedge \clk ) begin
        s63_val_n1 <= s62_val_n1;
    end
    always @(posedge \clk ) begin
        s63_val_n2 <= s62_val_n2;
    end
    always @(posedge \clk ) begin
        s63_val_n3 <= s62_val_n3;
    end
    always @(posedge \clk ) begin
        s63_val_n4 <= s62_val_n4;
    end
    always @(posedge \clk ) begin
        s63_val_n5 <= s62_val_n5;
    end
    always @(posedge \clk ) begin
        s63_val_n6 <= s62_val_n6;
    end
    always @(posedge \clk ) begin
        s63_val_n7 <= s62_val_n7;
    end
    always @(posedge \clk ) begin
        s63_val_n8 <= s62_val_n8;
    end
    always @(posedge \clk ) begin
        s63_val_n9 <= s62_val_n9;
    end
    always @(posedge \clk ) begin
        s63_val_n10 <= s62_val_n10;
    end
    always @(posedge \clk ) begin
        s63_val_n11 <= s62_val_n11;
    end
    always @(posedge \clk ) begin
        s63_val_n12 <= s62_val_n12;
    end
    always @(posedge \clk ) begin
        s63_val_n13 <= s62_val_n13;
    end
    always @(posedge \clk ) begin
        s63_val_n14 <= s62_val_n14;
    end
    always @(posedge \clk ) begin
        s63_val_n15 <= s62_val_n15;
    end
    always @(posedge \clk ) begin
        s63_val_n16 <= s62_val_n16;
    end
    always @(posedge \clk ) begin
        s63_val_n17 <= s62_val_n17;
    end
    always @(posedge \clk ) begin
        s63_val_n18 <= s62_val_n18;
    end
    always @(posedge \clk ) begin
        s63_val_n19 <= s62_val_n19;
    end
    always @(posedge \clk ) begin
        s63_val_n20 <= s62_val_n20;
    end
    always @(posedge \clk ) begin
        s63_val_n21 <= s62_val_n21;
    end
    always @(posedge \clk ) begin
        s63_val_n22 <= s62_val_n22;
    end
    always @(posedge \clk ) begin
        s63_val_n23 <= s62_val_n23;
    end
    always @(posedge \clk ) begin
        s63_val_n24 <= s62_val_n24;
    end
    always @(posedge \clk ) begin
        s63_val_n25 <= s62_val_n25;
    end
    always @(posedge \clk ) begin
        s63_val_n26 <= s62_val_n26;
    end
    always @(posedge \clk ) begin
        s63_val_n27 <= s62_val_n27;
    end
    always @(posedge \clk ) begin
        s63_val_n28 <= s62_val_n28;
    end
    always @(posedge \clk ) begin
        s63_val_n29 <= s62_val_n29;
    end
    always @(posedge \clk ) begin
        s63_val_n30 <= val_n30;
    end
    always @(posedge \clk ) begin
        \s64_val  <= \s63_val ;
    end
    always @(posedge \clk ) begin
        s64_val_n1 <= s63_val_n1;
    end
    always @(posedge \clk ) begin
        s64_val_n2 <= s63_val_n2;
    end
    always @(posedge \clk ) begin
        s64_val_n3 <= s63_val_n3;
    end
    always @(posedge \clk ) begin
        s64_val_n4 <= s63_val_n4;
    end
    always @(posedge \clk ) begin
        s64_val_n5 <= s63_val_n5;
    end
    always @(posedge \clk ) begin
        s64_val_n6 <= s63_val_n6;
    end
    always @(posedge \clk ) begin
        s64_val_n7 <= s63_val_n7;
    end
    always @(posedge \clk ) begin
        s64_val_n8 <= s63_val_n8;
    end
    always @(posedge \clk ) begin
        s64_val_n9 <= s63_val_n9;
    end
    always @(posedge \clk ) begin
        s64_val_n10 <= s63_val_n10;
    end
    always @(posedge \clk ) begin
        s64_val_n11 <= s63_val_n11;
    end
    always @(posedge \clk ) begin
        s64_val_n12 <= s63_val_n12;
    end
    always @(posedge \clk ) begin
        s64_val_n13 <= s63_val_n13;
    end
    always @(posedge \clk ) begin
        s64_val_n14 <= s63_val_n14;
    end
    always @(posedge \clk ) begin
        s64_val_n15 <= s63_val_n15;
    end
    always @(posedge \clk ) begin
        s64_val_n16 <= s63_val_n16;
    end
    always @(posedge \clk ) begin
        s64_val_n17 <= s63_val_n17;
    end
    always @(posedge \clk ) begin
        s64_val_n18 <= s63_val_n18;
    end
    always @(posedge \clk ) begin
        s64_val_n19 <= s63_val_n19;
    end
    always @(posedge \clk ) begin
        s64_val_n20 <= s63_val_n20;
    end
    always @(posedge \clk ) begin
        s64_val_n21 <= s63_val_n21;
    end
    always @(posedge \clk ) begin
        s64_val_n22 <= s63_val_n22;
    end
    always @(posedge \clk ) begin
        s64_val_n23 <= s63_val_n23;
    end
    always @(posedge \clk ) begin
        s64_val_n24 <= s63_val_n24;
    end
    always @(posedge \clk ) begin
        s64_val_n25 <= s63_val_n25;
    end
    always @(posedge \clk ) begin
        s64_val_n26 <= s63_val_n26;
    end
    always @(posedge \clk ) begin
        s64_val_n27 <= s63_val_n27;
    end
    always @(posedge \clk ) begin
        s64_val_n28 <= s63_val_n28;
    end
    always @(posedge \clk ) begin
        s64_val_n29 <= s63_val_n29;
    end
    always @(posedge \clk ) begin
        s64_val_n30 <= s63_val_n30;
    end
    always @(posedge \clk ) begin
        \s65_val  <= \s64_val ;
    end
    always @(posedge \clk ) begin
        s65_val_n1 <= s64_val_n1;
    end
    always @(posedge \clk ) begin
        s65_val_n2 <= s64_val_n2;
    end
    always @(posedge \clk ) begin
        s65_val_n3 <= s64_val_n3;
    end
    always @(posedge \clk ) begin
        s65_val_n4 <= s64_val_n4;
    end
    always @(posedge \clk ) begin
        s65_val_n5 <= s64_val_n5;
    end
    always @(posedge \clk ) begin
        s65_val_n6 <= s64_val_n6;
    end
    always @(posedge \clk ) begin
        s65_val_n7 <= s64_val_n7;
    end
    always @(posedge \clk ) begin
        s65_val_n8 <= s64_val_n8;
    end
    always @(posedge \clk ) begin
        s65_val_n9 <= s64_val_n9;
    end
    always @(posedge \clk ) begin
        s65_val_n10 <= s64_val_n10;
    end
    always @(posedge \clk ) begin
        s65_val_n11 <= s64_val_n11;
    end
    always @(posedge \clk ) begin
        s65_val_n12 <= s64_val_n12;
    end
    always @(posedge \clk ) begin
        s65_val_n13 <= s64_val_n13;
    end
    always @(posedge \clk ) begin
        s65_val_n14 <= s64_val_n14;
    end
    always @(posedge \clk ) begin
        s65_val_n15 <= s64_val_n15;
    end
    always @(posedge \clk ) begin
        s65_val_n16 <= s64_val_n16;
    end
    always @(posedge \clk ) begin
        s65_val_n17 <= s64_val_n17;
    end
    always @(posedge \clk ) begin
        s65_val_n18 <= s64_val_n18;
    end
    always @(posedge \clk ) begin
        s65_val_n19 <= s64_val_n19;
    end
    always @(posedge \clk ) begin
        s65_val_n20 <= s64_val_n20;
    end
    always @(posedge \clk ) begin
        s65_val_n21 <= s64_val_n21;
    end
    always @(posedge \clk ) begin
        s65_val_n22 <= s64_val_n22;
    end
    always @(posedge \clk ) begin
        s65_val_n23 <= s64_val_n23;
    end
    always @(posedge \clk ) begin
        s65_val_n24 <= s64_val_n24;
    end
    always @(posedge \clk ) begin
        s65_val_n25 <= s64_val_n25;
    end
    always @(posedge \clk ) begin
        s65_val_n26 <= s64_val_n26;
    end
    always @(posedge \clk ) begin
        s65_val_n27 <= s64_val_n27;
    end
    always @(posedge \clk ) begin
        s65_val_n28 <= s64_val_n28;
    end
    always @(posedge \clk ) begin
        s65_val_n29 <= s64_val_n29;
    end
    always @(posedge \clk ) begin
        s65_val_n30 <= s64_val_n30;
    end
    always @(posedge \clk ) begin
        s65_val_n31 <= val_n31;
    end
    always @(posedge \clk ) begin
        \s66_val  <= \s65_val ;
    end
    always @(posedge \clk ) begin
        s66_val_n1 <= s65_val_n1;
    end
    always @(posedge \clk ) begin
        s66_val_n2 <= s65_val_n2;
    end
    always @(posedge \clk ) begin
        s66_val_n3 <= s65_val_n3;
    end
    always @(posedge \clk ) begin
        s66_val_n4 <= s65_val_n4;
    end
    always @(posedge \clk ) begin
        s66_val_n5 <= s65_val_n5;
    end
    always @(posedge \clk ) begin
        s66_val_n6 <= s65_val_n6;
    end
    always @(posedge \clk ) begin
        s66_val_n7 <= s65_val_n7;
    end
    always @(posedge \clk ) begin
        s66_val_n8 <= s65_val_n8;
    end
    always @(posedge \clk ) begin
        s66_val_n9 <= s65_val_n9;
    end
    always @(posedge \clk ) begin
        s66_val_n10 <= s65_val_n10;
    end
    always @(posedge \clk ) begin
        s66_val_n11 <= s65_val_n11;
    end
    always @(posedge \clk ) begin
        s66_val_n12 <= s65_val_n12;
    end
    always @(posedge \clk ) begin
        s66_val_n13 <= s65_val_n13;
    end
    always @(posedge \clk ) begin
        s66_val_n14 <= s65_val_n14;
    end
    always @(posedge \clk ) begin
        s66_val_n15 <= s65_val_n15;
    end
    always @(posedge \clk ) begin
        s66_val_n16 <= s65_val_n16;
    end
    always @(posedge \clk ) begin
        s66_val_n17 <= s65_val_n17;
    end
    always @(posedge \clk ) begin
        s66_val_n18 <= s65_val_n18;
    end
    always @(posedge \clk ) begin
        s66_val_n19 <= s65_val_n19;
    end
    always @(posedge \clk ) begin
        s66_val_n20 <= s65_val_n20;
    end
    always @(posedge \clk ) begin
        s66_val_n21 <= s65_val_n21;
    end
    always @(posedge \clk ) begin
        s66_val_n22 <= s65_val_n22;
    end
    always @(posedge \clk ) begin
        s66_val_n23 <= s65_val_n23;
    end
    always @(posedge \clk ) begin
        s66_val_n24 <= s65_val_n24;
    end
    always @(posedge \clk ) begin
        s66_val_n25 <= s65_val_n25;
    end
    always @(posedge \clk ) begin
        s66_val_n26 <= s65_val_n26;
    end
    always @(posedge \clk ) begin
        s66_val_n27 <= s65_val_n27;
    end
    always @(posedge \clk ) begin
        s66_val_n28 <= s65_val_n28;
    end
    always @(posedge \clk ) begin
        s66_val_n29 <= s65_val_n29;
    end
    always @(posedge \clk ) begin
        s66_val_n30 <= s65_val_n30;
    end
    always @(posedge \clk ) begin
        s66_val_n31 <= s65_val_n31;
    end
    always @(posedge \clk ) begin
        \s67_val  <= \s66_val ;
    end
    always @(posedge \clk ) begin
        s67_val_n1 <= s66_val_n1;
    end
    always @(posedge \clk ) begin
        s67_val_n2 <= s66_val_n2;
    end
    always @(posedge \clk ) begin
        s67_val_n3 <= s66_val_n3;
    end
    always @(posedge \clk ) begin
        s67_val_n4 <= s66_val_n4;
    end
    always @(posedge \clk ) begin
        s67_val_n5 <= s66_val_n5;
    end
    always @(posedge \clk ) begin
        s67_val_n6 <= s66_val_n6;
    end
    always @(posedge \clk ) begin
        s67_val_n7 <= s66_val_n7;
    end
    always @(posedge \clk ) begin
        s67_val_n8 <= s66_val_n8;
    end
    always @(posedge \clk ) begin
        s67_val_n9 <= s66_val_n9;
    end
    always @(posedge \clk ) begin
        s67_val_n10 <= s66_val_n10;
    end
    always @(posedge \clk ) begin
        s67_val_n11 <= s66_val_n11;
    end
    always @(posedge \clk ) begin
        s67_val_n12 <= s66_val_n12;
    end
    always @(posedge \clk ) begin
        s67_val_n13 <= s66_val_n13;
    end
    always @(posedge \clk ) begin
        s67_val_n14 <= s66_val_n14;
    end
    always @(posedge \clk ) begin
        s67_val_n15 <= s66_val_n15;
    end
    always @(posedge \clk ) begin
        s67_val_n16 <= s66_val_n16;
    end
    always @(posedge \clk ) begin
        s67_val_n17 <= s66_val_n17;
    end
    always @(posedge \clk ) begin
        s67_val_n18 <= s66_val_n18;
    end
    always @(posedge \clk ) begin
        s67_val_n19 <= s66_val_n19;
    end
    always @(posedge \clk ) begin
        s67_val_n20 <= s66_val_n20;
    end
    always @(posedge \clk ) begin
        s67_val_n21 <= s66_val_n21;
    end
    always @(posedge \clk ) begin
        s67_val_n22 <= s66_val_n22;
    end
    always @(posedge \clk ) begin
        s67_val_n23 <= s66_val_n23;
    end
    always @(posedge \clk ) begin
        s67_val_n24 <= s66_val_n24;
    end
    always @(posedge \clk ) begin
        s67_val_n25 <= s66_val_n25;
    end
    always @(posedge \clk ) begin
        s67_val_n26 <= s66_val_n26;
    end
    always @(posedge \clk ) begin
        s67_val_n27 <= s66_val_n27;
    end
    always @(posedge \clk ) begin
        s67_val_n28 <= s66_val_n28;
    end
    always @(posedge \clk ) begin
        s67_val_n29 <= s66_val_n29;
    end
    always @(posedge \clk ) begin
        s67_val_n30 <= s66_val_n30;
    end
    always @(posedge \clk ) begin
        s67_val_n31 <= s66_val_n31;
    end
    always @(posedge \clk ) begin
        s67_val_n32 <= val_n32;
    end
    always @(posedge \clk ) begin
        \s68_val  <= \s67_val ;
    end
    always @(posedge \clk ) begin
        s68_val_n1 <= s67_val_n1;
    end
    always @(posedge \clk ) begin
        s68_val_n2 <= s67_val_n2;
    end
    always @(posedge \clk ) begin
        s68_val_n3 <= s67_val_n3;
    end
    always @(posedge \clk ) begin
        s68_val_n4 <= s67_val_n4;
    end
    always @(posedge \clk ) begin
        s68_val_n5 <= s67_val_n5;
    end
    always @(posedge \clk ) begin
        s68_val_n6 <= s67_val_n6;
    end
    always @(posedge \clk ) begin
        s68_val_n7 <= s67_val_n7;
    end
    always @(posedge \clk ) begin
        s68_val_n8 <= s67_val_n8;
    end
    always @(posedge \clk ) begin
        s68_val_n9 <= s67_val_n9;
    end
    always @(posedge \clk ) begin
        s68_val_n10 <= s67_val_n10;
    end
    always @(posedge \clk ) begin
        s68_val_n11 <= s67_val_n11;
    end
    always @(posedge \clk ) begin
        s68_val_n12 <= s67_val_n12;
    end
    always @(posedge \clk ) begin
        s68_val_n13 <= s67_val_n13;
    end
    always @(posedge \clk ) begin
        s68_val_n14 <= s67_val_n14;
    end
    always @(posedge \clk ) begin
        s68_val_n15 <= s67_val_n15;
    end
    always @(posedge \clk ) begin
        s68_val_n16 <= s67_val_n16;
    end
    always @(posedge \clk ) begin
        s68_val_n17 <= s67_val_n17;
    end
    always @(posedge \clk ) begin
        s68_val_n18 <= s67_val_n18;
    end
    always @(posedge \clk ) begin
        s68_val_n19 <= s67_val_n19;
    end
    always @(posedge \clk ) begin
        s68_val_n20 <= s67_val_n20;
    end
    always @(posedge \clk ) begin
        s68_val_n21 <= s67_val_n21;
    end
    always @(posedge \clk ) begin
        s68_val_n22 <= s67_val_n22;
    end
    always @(posedge \clk ) begin
        s68_val_n23 <= s67_val_n23;
    end
    always @(posedge \clk ) begin
        s68_val_n24 <= s67_val_n24;
    end
    always @(posedge \clk ) begin
        s68_val_n25 <= s67_val_n25;
    end
    always @(posedge \clk ) begin
        s68_val_n26 <= s67_val_n26;
    end
    always @(posedge \clk ) begin
        s68_val_n27 <= s67_val_n27;
    end
    always @(posedge \clk ) begin
        s68_val_n28 <= s67_val_n28;
    end
    always @(posedge \clk ) begin
        s68_val_n29 <= s67_val_n29;
    end
    always @(posedge \clk ) begin
        s68_val_n30 <= s67_val_n30;
    end
    always @(posedge \clk ) begin
        s68_val_n31 <= s67_val_n31;
    end
    always @(posedge \clk ) begin
        s68_val_n32 <= s67_val_n32;
    end
    always @(posedge \clk ) begin
        \s69_val  <= \s68_val ;
    end
    always @(posedge \clk ) begin
        s69_val_n1 <= s68_val_n1;
    end
    always @(posedge \clk ) begin
        s69_val_n2 <= s68_val_n2;
    end
    always @(posedge \clk ) begin
        s69_val_n3 <= s68_val_n3;
    end
    always @(posedge \clk ) begin
        s69_val_n4 <= s68_val_n4;
    end
    always @(posedge \clk ) begin
        s69_val_n5 <= s68_val_n5;
    end
    always @(posedge \clk ) begin
        s69_val_n6 <= s68_val_n6;
    end
    always @(posedge \clk ) begin
        s69_val_n7 <= s68_val_n7;
    end
    always @(posedge \clk ) begin
        s69_val_n8 <= s68_val_n8;
    end
    always @(posedge \clk ) begin
        s69_val_n9 <= s68_val_n9;
    end
    always @(posedge \clk ) begin
        s69_val_n10 <= s68_val_n10;
    end
    always @(posedge \clk ) begin
        s69_val_n11 <= s68_val_n11;
    end
    always @(posedge \clk ) begin
        s69_val_n12 <= s68_val_n12;
    end
    always @(posedge \clk ) begin
        s69_val_n13 <= s68_val_n13;
    end
    always @(posedge \clk ) begin
        s69_val_n14 <= s68_val_n14;
    end
    always @(posedge \clk ) begin
        s69_val_n15 <= s68_val_n15;
    end
    always @(posedge \clk ) begin
        s69_val_n16 <= s68_val_n16;
    end
    always @(posedge \clk ) begin
        s69_val_n17 <= s68_val_n17;
    end
    always @(posedge \clk ) begin
        s69_val_n18 <= s68_val_n18;
    end
    always @(posedge \clk ) begin
        s69_val_n19 <= s68_val_n19;
    end
    always @(posedge \clk ) begin
        s69_val_n20 <= s68_val_n20;
    end
    always @(posedge \clk ) begin
        s69_val_n21 <= s68_val_n21;
    end
    always @(posedge \clk ) begin
        s69_val_n22 <= s68_val_n22;
    end
    always @(posedge \clk ) begin
        s69_val_n23 <= s68_val_n23;
    end
    always @(posedge \clk ) begin
        s69_val_n24 <= s68_val_n24;
    end
    always @(posedge \clk ) begin
        s69_val_n25 <= s68_val_n25;
    end
    always @(posedge \clk ) begin
        s69_val_n26 <= s68_val_n26;
    end
    always @(posedge \clk ) begin
        s69_val_n27 <= s68_val_n27;
    end
    always @(posedge \clk ) begin
        s69_val_n28 <= s68_val_n28;
    end
    always @(posedge \clk ) begin
        s69_val_n29 <= s68_val_n29;
    end
    always @(posedge \clk ) begin
        s69_val_n30 <= s68_val_n30;
    end
    always @(posedge \clk ) begin
        s69_val_n31 <= s68_val_n31;
    end
    always @(posedge \clk ) begin
        s69_val_n32 <= s68_val_n32;
    end
    always @(posedge \clk ) begin
        s69_val_n33 <= val_n33;
    end
    always @(posedge \clk ) begin
        \s70_val  <= \s69_val ;
    end
    always @(posedge \clk ) begin
        s70_val_n1 <= s69_val_n1;
    end
    always @(posedge \clk ) begin
        s70_val_n2 <= s69_val_n2;
    end
    always @(posedge \clk ) begin
        s70_val_n3 <= s69_val_n3;
    end
    always @(posedge \clk ) begin
        s70_val_n4 <= s69_val_n4;
    end
    always @(posedge \clk ) begin
        s70_val_n5 <= s69_val_n5;
    end
    always @(posedge \clk ) begin
        s70_val_n6 <= s69_val_n6;
    end
    always @(posedge \clk ) begin
        s70_val_n7 <= s69_val_n7;
    end
    always @(posedge \clk ) begin
        s70_val_n8 <= s69_val_n8;
    end
    always @(posedge \clk ) begin
        s70_val_n9 <= s69_val_n9;
    end
    always @(posedge \clk ) begin
        s70_val_n10 <= s69_val_n10;
    end
    always @(posedge \clk ) begin
        s70_val_n11 <= s69_val_n11;
    end
    always @(posedge \clk ) begin
        s70_val_n12 <= s69_val_n12;
    end
    always @(posedge \clk ) begin
        s70_val_n13 <= s69_val_n13;
    end
    always @(posedge \clk ) begin
        s70_val_n14 <= s69_val_n14;
    end
    always @(posedge \clk ) begin
        s70_val_n15 <= s69_val_n15;
    end
    always @(posedge \clk ) begin
        s70_val_n16 <= s69_val_n16;
    end
    always @(posedge \clk ) begin
        s70_val_n17 <= s69_val_n17;
    end
    always @(posedge \clk ) begin
        s70_val_n18 <= s69_val_n18;
    end
    always @(posedge \clk ) begin
        s70_val_n19 <= s69_val_n19;
    end
    always @(posedge \clk ) begin
        s70_val_n20 <= s69_val_n20;
    end
    always @(posedge \clk ) begin
        s70_val_n21 <= s69_val_n21;
    end
    always @(posedge \clk ) begin
        s70_val_n22 <= s69_val_n22;
    end
    always @(posedge \clk ) begin
        s70_val_n23 <= s69_val_n23;
    end
    always @(posedge \clk ) begin
        s70_val_n24 <= s69_val_n24;
    end
    always @(posedge \clk ) begin
        s70_val_n25 <= s69_val_n25;
    end
    always @(posedge \clk ) begin
        s70_val_n26 <= s69_val_n26;
    end
    always @(posedge \clk ) begin
        s70_val_n27 <= s69_val_n27;
    end
    always @(posedge \clk ) begin
        s70_val_n28 <= s69_val_n28;
    end
    always @(posedge \clk ) begin
        s70_val_n29 <= s69_val_n29;
    end
    always @(posedge \clk ) begin
        s70_val_n30 <= s69_val_n30;
    end
    always @(posedge \clk ) begin
        s70_val_n31 <= s69_val_n31;
    end
    always @(posedge \clk ) begin
        s70_val_n32 <= s69_val_n32;
    end
    always @(posedge \clk ) begin
        s70_val_n33 <= s69_val_n33;
    end
    always @(posedge \clk ) begin
        \s71_val  <= \s70_val ;
    end
    always @(posedge \clk ) begin
        s71_val_n1 <= s70_val_n1;
    end
    always @(posedge \clk ) begin
        s71_val_n2 <= s70_val_n2;
    end
    always @(posedge \clk ) begin
        s71_val_n3 <= s70_val_n3;
    end
    always @(posedge \clk ) begin
        s71_val_n4 <= s70_val_n4;
    end
    always @(posedge \clk ) begin
        s71_val_n5 <= s70_val_n5;
    end
    always @(posedge \clk ) begin
        s71_val_n6 <= s70_val_n6;
    end
    always @(posedge \clk ) begin
        s71_val_n7 <= s70_val_n7;
    end
    always @(posedge \clk ) begin
        s71_val_n8 <= s70_val_n8;
    end
    always @(posedge \clk ) begin
        s71_val_n9 <= s70_val_n9;
    end
    always @(posedge \clk ) begin
        s71_val_n10 <= s70_val_n10;
    end
    always @(posedge \clk ) begin
        s71_val_n11 <= s70_val_n11;
    end
    always @(posedge \clk ) begin
        s71_val_n12 <= s70_val_n12;
    end
    always @(posedge \clk ) begin
        s71_val_n13 <= s70_val_n13;
    end
    always @(posedge \clk ) begin
        s71_val_n14 <= s70_val_n14;
    end
    always @(posedge \clk ) begin
        s71_val_n15 <= s70_val_n15;
    end
    always @(posedge \clk ) begin
        s71_val_n16 <= s70_val_n16;
    end
    always @(posedge \clk ) begin
        s71_val_n17 <= s70_val_n17;
    end
    always @(posedge \clk ) begin
        s71_val_n18 <= s70_val_n18;
    end
    always @(posedge \clk ) begin
        s71_val_n19 <= s70_val_n19;
    end
    always @(posedge \clk ) begin
        s71_val_n20 <= s70_val_n20;
    end
    always @(posedge \clk ) begin
        s71_val_n21 <= s70_val_n21;
    end
    always @(posedge \clk ) begin
        s71_val_n22 <= s70_val_n22;
    end
    always @(posedge \clk ) begin
        s71_val_n23 <= s70_val_n23;
    end
    always @(posedge \clk ) begin
        s71_val_n24 <= s70_val_n24;
    end
    always @(posedge \clk ) begin
        s71_val_n25 <= s70_val_n25;
    end
    always @(posedge \clk ) begin
        s71_val_n26 <= s70_val_n26;
    end
    always @(posedge \clk ) begin
        s71_val_n27 <= s70_val_n27;
    end
    always @(posedge \clk ) begin
        s71_val_n28 <= s70_val_n28;
    end
    always @(posedge \clk ) begin
        s71_val_n29 <= s70_val_n29;
    end
    always @(posedge \clk ) begin
        s71_val_n30 <= s70_val_n30;
    end
    always @(posedge \clk ) begin
        s71_val_n31 <= s70_val_n31;
    end
    always @(posedge \clk ) begin
        s71_val_n32 <= s70_val_n32;
    end
    always @(posedge \clk ) begin
        s71_val_n33 <= s70_val_n33;
    end
    always @(posedge \clk ) begin
        s71_val_n34 <= val_n34;
    end
    always @(posedge \clk ) begin
        \s72_val  <= \s71_val ;
    end
    always @(posedge \clk ) begin
        s72_val_n1 <= s71_val_n1;
    end
    always @(posedge \clk ) begin
        s72_val_n2 <= s71_val_n2;
    end
    always @(posedge \clk ) begin
        s72_val_n3 <= s71_val_n3;
    end
    always @(posedge \clk ) begin
        s72_val_n4 <= s71_val_n4;
    end
    always @(posedge \clk ) begin
        s72_val_n5 <= s71_val_n5;
    end
    always @(posedge \clk ) begin
        s72_val_n6 <= s71_val_n6;
    end
    always @(posedge \clk ) begin
        s72_val_n7 <= s71_val_n7;
    end
    always @(posedge \clk ) begin
        s72_val_n8 <= s71_val_n8;
    end
    always @(posedge \clk ) begin
        s72_val_n9 <= s71_val_n9;
    end
    always @(posedge \clk ) begin
        s72_val_n10 <= s71_val_n10;
    end
    always @(posedge \clk ) begin
        s72_val_n11 <= s71_val_n11;
    end
    always @(posedge \clk ) begin
        s72_val_n12 <= s71_val_n12;
    end
    always @(posedge \clk ) begin
        s72_val_n13 <= s71_val_n13;
    end
    always @(posedge \clk ) begin
        s72_val_n14 <= s71_val_n14;
    end
    always @(posedge \clk ) begin
        s72_val_n15 <= s71_val_n15;
    end
    always @(posedge \clk ) begin
        s72_val_n16 <= s71_val_n16;
    end
    always @(posedge \clk ) begin
        s72_val_n17 <= s71_val_n17;
    end
    always @(posedge \clk ) begin
        s72_val_n18 <= s71_val_n18;
    end
    always @(posedge \clk ) begin
        s72_val_n19 <= s71_val_n19;
    end
    always @(posedge \clk ) begin
        s72_val_n20 <= s71_val_n20;
    end
    always @(posedge \clk ) begin
        s72_val_n21 <= s71_val_n21;
    end
    always @(posedge \clk ) begin
        s72_val_n22 <= s71_val_n22;
    end
    always @(posedge \clk ) begin
        s72_val_n23 <= s71_val_n23;
    end
    always @(posedge \clk ) begin
        s72_val_n24 <= s71_val_n24;
    end
    always @(posedge \clk ) begin
        s72_val_n25 <= s71_val_n25;
    end
    always @(posedge \clk ) begin
        s72_val_n26 <= s71_val_n26;
    end
    always @(posedge \clk ) begin
        s72_val_n27 <= s71_val_n27;
    end
    always @(posedge \clk ) begin
        s72_val_n28 <= s71_val_n28;
    end
    always @(posedge \clk ) begin
        s72_val_n29 <= s71_val_n29;
    end
    always @(posedge \clk ) begin
        s72_val_n30 <= s71_val_n30;
    end
    always @(posedge \clk ) begin
        s72_val_n31 <= s71_val_n31;
    end
    always @(posedge \clk ) begin
        s72_val_n32 <= s71_val_n32;
    end
    always @(posedge \clk ) begin
        s72_val_n33 <= s71_val_n33;
    end
    always @(posedge \clk ) begin
        s72_val_n34 <= s71_val_n34;
    end
    always @(posedge \clk ) begin
        \s73_val  <= \s72_val ;
    end
    always @(posedge \clk ) begin
        s73_val_n1 <= s72_val_n1;
    end
    always @(posedge \clk ) begin
        s73_val_n2 <= s72_val_n2;
    end
    always @(posedge \clk ) begin
        s73_val_n3 <= s72_val_n3;
    end
    always @(posedge \clk ) begin
        s73_val_n4 <= s72_val_n4;
    end
    always @(posedge \clk ) begin
        s73_val_n5 <= s72_val_n5;
    end
    always @(posedge \clk ) begin
        s73_val_n6 <= s72_val_n6;
    end
    always @(posedge \clk ) begin
        s73_val_n7 <= s72_val_n7;
    end
    always @(posedge \clk ) begin
        s73_val_n8 <= s72_val_n8;
    end
    always @(posedge \clk ) begin
        s73_val_n9 <= s72_val_n9;
    end
    always @(posedge \clk ) begin
        s73_val_n10 <= s72_val_n10;
    end
    always @(posedge \clk ) begin
        s73_val_n11 <= s72_val_n11;
    end
    always @(posedge \clk ) begin
        s73_val_n12 <= s72_val_n12;
    end
    always @(posedge \clk ) begin
        s73_val_n13 <= s72_val_n13;
    end
    always @(posedge \clk ) begin
        s73_val_n14 <= s72_val_n14;
    end
    always @(posedge \clk ) begin
        s73_val_n15 <= s72_val_n15;
    end
    always @(posedge \clk ) begin
        s73_val_n16 <= s72_val_n16;
    end
    always @(posedge \clk ) begin
        s73_val_n17 <= s72_val_n17;
    end
    always @(posedge \clk ) begin
        s73_val_n18 <= s72_val_n18;
    end
    always @(posedge \clk ) begin
        s73_val_n19 <= s72_val_n19;
    end
    always @(posedge \clk ) begin
        s73_val_n20 <= s72_val_n20;
    end
    always @(posedge \clk ) begin
        s73_val_n21 <= s72_val_n21;
    end
    always @(posedge \clk ) begin
        s73_val_n22 <= s72_val_n22;
    end
    always @(posedge \clk ) begin
        s73_val_n23 <= s72_val_n23;
    end
    always @(posedge \clk ) begin
        s73_val_n24 <= s72_val_n24;
    end
    always @(posedge \clk ) begin
        s73_val_n25 <= s72_val_n25;
    end
    always @(posedge \clk ) begin
        s73_val_n26 <= s72_val_n26;
    end
    always @(posedge \clk ) begin
        s73_val_n27 <= s72_val_n27;
    end
    always @(posedge \clk ) begin
        s73_val_n28 <= s72_val_n28;
    end
    always @(posedge \clk ) begin
        s73_val_n29 <= s72_val_n29;
    end
    always @(posedge \clk ) begin
        s73_val_n30 <= s72_val_n30;
    end
    always @(posedge \clk ) begin
        s73_val_n31 <= s72_val_n31;
    end
    always @(posedge \clk ) begin
        s73_val_n32 <= s72_val_n32;
    end
    always @(posedge \clk ) begin
        s73_val_n33 <= s72_val_n33;
    end
    always @(posedge \clk ) begin
        s73_val_n34 <= s72_val_n34;
    end
    always @(posedge \clk ) begin
        s73_val_n35 <= val_n35;
    end
    always @(posedge \clk ) begin
        \s74_val  <= \s73_val ;
    end
    always @(posedge \clk ) begin
        s74_val_n1 <= s73_val_n1;
    end
    always @(posedge \clk ) begin
        s74_val_n2 <= s73_val_n2;
    end
    always @(posedge \clk ) begin
        s74_val_n3 <= s73_val_n3;
    end
    always @(posedge \clk ) begin
        s74_val_n4 <= s73_val_n4;
    end
    always @(posedge \clk ) begin
        s74_val_n5 <= s73_val_n5;
    end
    always @(posedge \clk ) begin
        s74_val_n6 <= s73_val_n6;
    end
    always @(posedge \clk ) begin
        s74_val_n7 <= s73_val_n7;
    end
    always @(posedge \clk ) begin
        s74_val_n8 <= s73_val_n8;
    end
    always @(posedge \clk ) begin
        s74_val_n9 <= s73_val_n9;
    end
    always @(posedge \clk ) begin
        s74_val_n10 <= s73_val_n10;
    end
    always @(posedge \clk ) begin
        s74_val_n11 <= s73_val_n11;
    end
    always @(posedge \clk ) begin
        s74_val_n12 <= s73_val_n12;
    end
    always @(posedge \clk ) begin
        s74_val_n13 <= s73_val_n13;
    end
    always @(posedge \clk ) begin
        s74_val_n14 <= s73_val_n14;
    end
    always @(posedge \clk ) begin
        s74_val_n15 <= s73_val_n15;
    end
    always @(posedge \clk ) begin
        s74_val_n16 <= s73_val_n16;
    end
    always @(posedge \clk ) begin
        s74_val_n17 <= s73_val_n17;
    end
    always @(posedge \clk ) begin
        s74_val_n18 <= s73_val_n18;
    end
    always @(posedge \clk ) begin
        s74_val_n19 <= s73_val_n19;
    end
    always @(posedge \clk ) begin
        s74_val_n20 <= s73_val_n20;
    end
    always @(posedge \clk ) begin
        s74_val_n21 <= s73_val_n21;
    end
    always @(posedge \clk ) begin
        s74_val_n22 <= s73_val_n22;
    end
    always @(posedge \clk ) begin
        s74_val_n23 <= s73_val_n23;
    end
    always @(posedge \clk ) begin
        s74_val_n24 <= s73_val_n24;
    end
    always @(posedge \clk ) begin
        s74_val_n25 <= s73_val_n25;
    end
    always @(posedge \clk ) begin
        s74_val_n26 <= s73_val_n26;
    end
    always @(posedge \clk ) begin
        s74_val_n27 <= s73_val_n27;
    end
    always @(posedge \clk ) begin
        s74_val_n28 <= s73_val_n28;
    end
    always @(posedge \clk ) begin
        s74_val_n29 <= s73_val_n29;
    end
    always @(posedge \clk ) begin
        s74_val_n30 <= s73_val_n30;
    end
    always @(posedge \clk ) begin
        s74_val_n31 <= s73_val_n31;
    end
    always @(posedge \clk ) begin
        s74_val_n32 <= s73_val_n32;
    end
    always @(posedge \clk ) begin
        s74_val_n33 <= s73_val_n33;
    end
    always @(posedge \clk ) begin
        s74_val_n34 <= s73_val_n34;
    end
    always @(posedge \clk ) begin
        s74_val_n35 <= s73_val_n35;
    end
    always @(posedge \clk ) begin
        \s75_val  <= \s74_val ;
    end
    always @(posedge \clk ) begin
        s75_val_n1 <= s74_val_n1;
    end
    always @(posedge \clk ) begin
        s75_val_n2 <= s74_val_n2;
    end
    always @(posedge \clk ) begin
        s75_val_n3 <= s74_val_n3;
    end
    always @(posedge \clk ) begin
        s75_val_n4 <= s74_val_n4;
    end
    always @(posedge \clk ) begin
        s75_val_n5 <= s74_val_n5;
    end
    always @(posedge \clk ) begin
        s75_val_n6 <= s74_val_n6;
    end
    always @(posedge \clk ) begin
        s75_val_n7 <= s74_val_n7;
    end
    always @(posedge \clk ) begin
        s75_val_n8 <= s74_val_n8;
    end
    always @(posedge \clk ) begin
        s75_val_n9 <= s74_val_n9;
    end
    always @(posedge \clk ) begin
        s75_val_n10 <= s74_val_n10;
    end
    always @(posedge \clk ) begin
        s75_val_n11 <= s74_val_n11;
    end
    always @(posedge \clk ) begin
        s75_val_n12 <= s74_val_n12;
    end
    always @(posedge \clk ) begin
        s75_val_n13 <= s74_val_n13;
    end
    always @(posedge \clk ) begin
        s75_val_n14 <= s74_val_n14;
    end
    always @(posedge \clk ) begin
        s75_val_n15 <= s74_val_n15;
    end
    always @(posedge \clk ) begin
        s75_val_n16 <= s74_val_n16;
    end
    always @(posedge \clk ) begin
        s75_val_n17 <= s74_val_n17;
    end
    always @(posedge \clk ) begin
        s75_val_n18 <= s74_val_n18;
    end
    always @(posedge \clk ) begin
        s75_val_n19 <= s74_val_n19;
    end
    always @(posedge \clk ) begin
        s75_val_n20 <= s74_val_n20;
    end
    always @(posedge \clk ) begin
        s75_val_n21 <= s74_val_n21;
    end
    always @(posedge \clk ) begin
        s75_val_n22 <= s74_val_n22;
    end
    always @(posedge \clk ) begin
        s75_val_n23 <= s74_val_n23;
    end
    always @(posedge \clk ) begin
        s75_val_n24 <= s74_val_n24;
    end
    always @(posedge \clk ) begin
        s75_val_n25 <= s74_val_n25;
    end
    always @(posedge \clk ) begin
        s75_val_n26 <= s74_val_n26;
    end
    always @(posedge \clk ) begin
        s75_val_n27 <= s74_val_n27;
    end
    always @(posedge \clk ) begin
        s75_val_n28 <= s74_val_n28;
    end
    always @(posedge \clk ) begin
        s75_val_n29 <= s74_val_n29;
    end
    always @(posedge \clk ) begin
        s75_val_n30 <= s74_val_n30;
    end
    always @(posedge \clk ) begin
        s75_val_n31 <= s74_val_n31;
    end
    always @(posedge \clk ) begin
        s75_val_n32 <= s74_val_n32;
    end
    always @(posedge \clk ) begin
        s75_val_n33 <= s74_val_n33;
    end
    always @(posedge \clk ) begin
        s75_val_n34 <= s74_val_n34;
    end
    always @(posedge \clk ) begin
        s75_val_n35 <= s74_val_n35;
    end
    always @(posedge \clk ) begin
        s75_val_n36 <= val_n36;
    end
    always @(posedge \clk ) begin
        \s76_val  <= \s75_val ;
    end
    always @(posedge \clk ) begin
        s76_val_n1 <= s75_val_n1;
    end
    always @(posedge \clk ) begin
        s76_val_n2 <= s75_val_n2;
    end
    always @(posedge \clk ) begin
        s76_val_n3 <= s75_val_n3;
    end
    always @(posedge \clk ) begin
        s76_val_n4 <= s75_val_n4;
    end
    always @(posedge \clk ) begin
        s76_val_n5 <= s75_val_n5;
    end
    always @(posedge \clk ) begin
        s76_val_n6 <= s75_val_n6;
    end
    always @(posedge \clk ) begin
        s76_val_n7 <= s75_val_n7;
    end
    always @(posedge \clk ) begin
        s76_val_n8 <= s75_val_n8;
    end
    always @(posedge \clk ) begin
        s76_val_n9 <= s75_val_n9;
    end
    always @(posedge \clk ) begin
        s76_val_n10 <= s75_val_n10;
    end
    always @(posedge \clk ) begin
        s76_val_n11 <= s75_val_n11;
    end
    always @(posedge \clk ) begin
        s76_val_n12 <= s75_val_n12;
    end
    always @(posedge \clk ) begin
        s76_val_n13 <= s75_val_n13;
    end
    always @(posedge \clk ) begin
        s76_val_n14 <= s75_val_n14;
    end
    always @(posedge \clk ) begin
        s76_val_n15 <= s75_val_n15;
    end
    always @(posedge \clk ) begin
        s76_val_n16 <= s75_val_n16;
    end
    always @(posedge \clk ) begin
        s76_val_n17 <= s75_val_n17;
    end
    always @(posedge \clk ) begin
        s76_val_n18 <= s75_val_n18;
    end
    always @(posedge \clk ) begin
        s76_val_n19 <= s75_val_n19;
    end
    always @(posedge \clk ) begin
        s76_val_n20 <= s75_val_n20;
    end
    always @(posedge \clk ) begin
        s76_val_n21 <= s75_val_n21;
    end
    always @(posedge \clk ) begin
        s76_val_n22 <= s75_val_n22;
    end
    always @(posedge \clk ) begin
        s76_val_n23 <= s75_val_n23;
    end
    always @(posedge \clk ) begin
        s76_val_n24 <= s75_val_n24;
    end
    always @(posedge \clk ) begin
        s76_val_n25 <= s75_val_n25;
    end
    always @(posedge \clk ) begin
        s76_val_n26 <= s75_val_n26;
    end
    always @(posedge \clk ) begin
        s76_val_n27 <= s75_val_n27;
    end
    always @(posedge \clk ) begin
        s76_val_n28 <= s75_val_n28;
    end
    always @(posedge \clk ) begin
        s76_val_n29 <= s75_val_n29;
    end
    always @(posedge \clk ) begin
        s76_val_n30 <= s75_val_n30;
    end
    always @(posedge \clk ) begin
        s76_val_n31 <= s75_val_n31;
    end
    always @(posedge \clk ) begin
        s76_val_n32 <= s75_val_n32;
    end
    always @(posedge \clk ) begin
        s76_val_n33 <= s75_val_n33;
    end
    always @(posedge \clk ) begin
        s76_val_n34 <= s75_val_n34;
    end
    always @(posedge \clk ) begin
        s76_val_n35 <= s75_val_n35;
    end
    always @(posedge \clk ) begin
        s76_val_n36 <= s75_val_n36;
    end
    always @(posedge \clk ) begin
        \s77_val  <= \s76_val ;
    end
    always @(posedge \clk ) begin
        s77_val_n1 <= s76_val_n1;
    end
    always @(posedge \clk ) begin
        s77_val_n2 <= s76_val_n2;
    end
    always @(posedge \clk ) begin
        s77_val_n3 <= s76_val_n3;
    end
    always @(posedge \clk ) begin
        s77_val_n4 <= s76_val_n4;
    end
    always @(posedge \clk ) begin
        s77_val_n5 <= s76_val_n5;
    end
    always @(posedge \clk ) begin
        s77_val_n6 <= s76_val_n6;
    end
    always @(posedge \clk ) begin
        s77_val_n7 <= s76_val_n7;
    end
    always @(posedge \clk ) begin
        s77_val_n8 <= s76_val_n8;
    end
    always @(posedge \clk ) begin
        s77_val_n9 <= s76_val_n9;
    end
    always @(posedge \clk ) begin
        s77_val_n10 <= s76_val_n10;
    end
    always @(posedge \clk ) begin
        s77_val_n11 <= s76_val_n11;
    end
    always @(posedge \clk ) begin
        s77_val_n12 <= s76_val_n12;
    end
    always @(posedge \clk ) begin
        s77_val_n13 <= s76_val_n13;
    end
    always @(posedge \clk ) begin
        s77_val_n14 <= s76_val_n14;
    end
    always @(posedge \clk ) begin
        s77_val_n15 <= s76_val_n15;
    end
    always @(posedge \clk ) begin
        s77_val_n16 <= s76_val_n16;
    end
    always @(posedge \clk ) begin
        s77_val_n17 <= s76_val_n17;
    end
    always @(posedge \clk ) begin
        s77_val_n18 <= s76_val_n18;
    end
    always @(posedge \clk ) begin
        s77_val_n19 <= s76_val_n19;
    end
    always @(posedge \clk ) begin
        s77_val_n20 <= s76_val_n20;
    end
    always @(posedge \clk ) begin
        s77_val_n21 <= s76_val_n21;
    end
    always @(posedge \clk ) begin
        s77_val_n22 <= s76_val_n22;
    end
    always @(posedge \clk ) begin
        s77_val_n23 <= s76_val_n23;
    end
    always @(posedge \clk ) begin
        s77_val_n24 <= s76_val_n24;
    end
    always @(posedge \clk ) begin
        s77_val_n25 <= s76_val_n25;
    end
    always @(posedge \clk ) begin
        s77_val_n26 <= s76_val_n26;
    end
    always @(posedge \clk ) begin
        s77_val_n27 <= s76_val_n27;
    end
    always @(posedge \clk ) begin
        s77_val_n28 <= s76_val_n28;
    end
    always @(posedge \clk ) begin
        s77_val_n29 <= s76_val_n29;
    end
    always @(posedge \clk ) begin
        s77_val_n30 <= s76_val_n30;
    end
    always @(posedge \clk ) begin
        s77_val_n31 <= s76_val_n31;
    end
    always @(posedge \clk ) begin
        s77_val_n32 <= s76_val_n32;
    end
    always @(posedge \clk ) begin
        s77_val_n33 <= s76_val_n33;
    end
    always @(posedge \clk ) begin
        s77_val_n34 <= s76_val_n34;
    end
    always @(posedge \clk ) begin
        s77_val_n35 <= s76_val_n35;
    end
    always @(posedge \clk ) begin
        s77_val_n36 <= s76_val_n36;
    end
    always @(posedge \clk ) begin
        s77_val_n37 <= val_n37;
    end
    always @(posedge \clk ) begin
        \s78_val  <= \s77_val ;
    end
    always @(posedge \clk ) begin
        s78_val_n1 <= s77_val_n1;
    end
    always @(posedge \clk ) begin
        s78_val_n2 <= s77_val_n2;
    end
    always @(posedge \clk ) begin
        s78_val_n3 <= s77_val_n3;
    end
    always @(posedge \clk ) begin
        s78_val_n4 <= s77_val_n4;
    end
    always @(posedge \clk ) begin
        s78_val_n5 <= s77_val_n5;
    end
    always @(posedge \clk ) begin
        s78_val_n6 <= s77_val_n6;
    end
    always @(posedge \clk ) begin
        s78_val_n7 <= s77_val_n7;
    end
    always @(posedge \clk ) begin
        s78_val_n8 <= s77_val_n8;
    end
    always @(posedge \clk ) begin
        s78_val_n9 <= s77_val_n9;
    end
    always @(posedge \clk ) begin
        s78_val_n10 <= s77_val_n10;
    end
    always @(posedge \clk ) begin
        s78_val_n11 <= s77_val_n11;
    end
    always @(posedge \clk ) begin
        s78_val_n12 <= s77_val_n12;
    end
    always @(posedge \clk ) begin
        s78_val_n13 <= s77_val_n13;
    end
    always @(posedge \clk ) begin
        s78_val_n14 <= s77_val_n14;
    end
    always @(posedge \clk ) begin
        s78_val_n15 <= s77_val_n15;
    end
    always @(posedge \clk ) begin
        s78_val_n16 <= s77_val_n16;
    end
    always @(posedge \clk ) begin
        s78_val_n17 <= s77_val_n17;
    end
    always @(posedge \clk ) begin
        s78_val_n18 <= s77_val_n18;
    end
    always @(posedge \clk ) begin
        s78_val_n19 <= s77_val_n19;
    end
    always @(posedge \clk ) begin
        s78_val_n20 <= s77_val_n20;
    end
    always @(posedge \clk ) begin
        s78_val_n21 <= s77_val_n21;
    end
    always @(posedge \clk ) begin
        s78_val_n22 <= s77_val_n22;
    end
    always @(posedge \clk ) begin
        s78_val_n23 <= s77_val_n23;
    end
    always @(posedge \clk ) begin
        s78_val_n24 <= s77_val_n24;
    end
    always @(posedge \clk ) begin
        s78_val_n25 <= s77_val_n25;
    end
    always @(posedge \clk ) begin
        s78_val_n26 <= s77_val_n26;
    end
    always @(posedge \clk ) begin
        s78_val_n27 <= s77_val_n27;
    end
    always @(posedge \clk ) begin
        s78_val_n28 <= s77_val_n28;
    end
    always @(posedge \clk ) begin
        s78_val_n29 <= s77_val_n29;
    end
    always @(posedge \clk ) begin
        s78_val_n30 <= s77_val_n30;
    end
    always @(posedge \clk ) begin
        s78_val_n31 <= s77_val_n31;
    end
    always @(posedge \clk ) begin
        s78_val_n32 <= s77_val_n32;
    end
    always @(posedge \clk ) begin
        s78_val_n33 <= s77_val_n33;
    end
    always @(posedge \clk ) begin
        s78_val_n34 <= s77_val_n34;
    end
    always @(posedge \clk ) begin
        s78_val_n35 <= s77_val_n35;
    end
    always @(posedge \clk ) begin
        s78_val_n36 <= s77_val_n36;
    end
    always @(posedge \clk ) begin
        s78_val_n37 <= s77_val_n37;
    end
    always @(posedge \clk ) begin
        \s79_val  <= \s78_val ;
    end
    always @(posedge \clk ) begin
        s79_val_n1 <= s78_val_n1;
    end
    always @(posedge \clk ) begin
        s79_val_n2 <= s78_val_n2;
    end
    always @(posedge \clk ) begin
        s79_val_n3 <= s78_val_n3;
    end
    always @(posedge \clk ) begin
        s79_val_n4 <= s78_val_n4;
    end
    always @(posedge \clk ) begin
        s79_val_n5 <= s78_val_n5;
    end
    always @(posedge \clk ) begin
        s79_val_n6 <= s78_val_n6;
    end
    always @(posedge \clk ) begin
        s79_val_n7 <= s78_val_n7;
    end
    always @(posedge \clk ) begin
        s79_val_n8 <= s78_val_n8;
    end
    always @(posedge \clk ) begin
        s79_val_n9 <= s78_val_n9;
    end
    always @(posedge \clk ) begin
        s79_val_n10 <= s78_val_n10;
    end
    always @(posedge \clk ) begin
        s79_val_n11 <= s78_val_n11;
    end
    always @(posedge \clk ) begin
        s79_val_n12 <= s78_val_n12;
    end
    always @(posedge \clk ) begin
        s79_val_n13 <= s78_val_n13;
    end
    always @(posedge \clk ) begin
        s79_val_n14 <= s78_val_n14;
    end
    always @(posedge \clk ) begin
        s79_val_n15 <= s78_val_n15;
    end
    always @(posedge \clk ) begin
        s79_val_n16 <= s78_val_n16;
    end
    always @(posedge \clk ) begin
        s79_val_n17 <= s78_val_n17;
    end
    always @(posedge \clk ) begin
        s79_val_n18 <= s78_val_n18;
    end
    always @(posedge \clk ) begin
        s79_val_n19 <= s78_val_n19;
    end
    always @(posedge \clk ) begin
        s79_val_n20 <= s78_val_n20;
    end
    always @(posedge \clk ) begin
        s79_val_n21 <= s78_val_n21;
    end
    always @(posedge \clk ) begin
        s79_val_n22 <= s78_val_n22;
    end
    always @(posedge \clk ) begin
        s79_val_n23 <= s78_val_n23;
    end
    always @(posedge \clk ) begin
        s79_val_n24 <= s78_val_n24;
    end
    always @(posedge \clk ) begin
        s79_val_n25 <= s78_val_n25;
    end
    always @(posedge \clk ) begin
        s79_val_n26 <= s78_val_n26;
    end
    always @(posedge \clk ) begin
        s79_val_n27 <= s78_val_n27;
    end
    always @(posedge \clk ) begin
        s79_val_n28 <= s78_val_n28;
    end
    always @(posedge \clk ) begin
        s79_val_n29 <= s78_val_n29;
    end
    always @(posedge \clk ) begin
        s79_val_n30 <= s78_val_n30;
    end
    always @(posedge \clk ) begin
        s79_val_n31 <= s78_val_n31;
    end
    always @(posedge \clk ) begin
        s79_val_n32 <= s78_val_n32;
    end
    always @(posedge \clk ) begin
        s79_val_n33 <= s78_val_n33;
    end
    always @(posedge \clk ) begin
        s79_val_n34 <= s78_val_n34;
    end
    always @(posedge \clk ) begin
        s79_val_n35 <= s78_val_n35;
    end
    always @(posedge \clk ) begin
        s79_val_n36 <= s78_val_n36;
    end
    always @(posedge \clk ) begin
        s79_val_n37 <= s78_val_n37;
    end
    always @(posedge \clk ) begin
        s79_val_n38 <= val_n38;
    end
    always @(posedge \clk ) begin
        \s80_val  <= \s79_val ;
    end
    always @(posedge \clk ) begin
        s80_val_n1 <= s79_val_n1;
    end
    always @(posedge \clk ) begin
        s80_val_n2 <= s79_val_n2;
    end
    always @(posedge \clk ) begin
        s80_val_n3 <= s79_val_n3;
    end
    always @(posedge \clk ) begin
        s80_val_n4 <= s79_val_n4;
    end
    always @(posedge \clk ) begin
        s80_val_n5 <= s79_val_n5;
    end
    always @(posedge \clk ) begin
        s80_val_n6 <= s79_val_n6;
    end
    always @(posedge \clk ) begin
        s80_val_n7 <= s79_val_n7;
    end
    always @(posedge \clk ) begin
        s80_val_n8 <= s79_val_n8;
    end
    always @(posedge \clk ) begin
        s80_val_n9 <= s79_val_n9;
    end
    always @(posedge \clk ) begin
        s80_val_n10 <= s79_val_n10;
    end
    always @(posedge \clk ) begin
        s80_val_n11 <= s79_val_n11;
    end
    always @(posedge \clk ) begin
        s80_val_n12 <= s79_val_n12;
    end
    always @(posedge \clk ) begin
        s80_val_n13 <= s79_val_n13;
    end
    always @(posedge \clk ) begin
        s80_val_n14 <= s79_val_n14;
    end
    always @(posedge \clk ) begin
        s80_val_n15 <= s79_val_n15;
    end
    always @(posedge \clk ) begin
        s80_val_n16 <= s79_val_n16;
    end
    always @(posedge \clk ) begin
        s80_val_n17 <= s79_val_n17;
    end
    always @(posedge \clk ) begin
        s80_val_n18 <= s79_val_n18;
    end
    always @(posedge \clk ) begin
        s80_val_n19 <= s79_val_n19;
    end
    always @(posedge \clk ) begin
        s80_val_n20 <= s79_val_n20;
    end
    always @(posedge \clk ) begin
        s80_val_n21 <= s79_val_n21;
    end
    always @(posedge \clk ) begin
        s80_val_n22 <= s79_val_n22;
    end
    always @(posedge \clk ) begin
        s80_val_n23 <= s79_val_n23;
    end
    always @(posedge \clk ) begin
        s80_val_n24 <= s79_val_n24;
    end
    always @(posedge \clk ) begin
        s80_val_n25 <= s79_val_n25;
    end
    always @(posedge \clk ) begin
        s80_val_n26 <= s79_val_n26;
    end
    always @(posedge \clk ) begin
        s80_val_n27 <= s79_val_n27;
    end
    always @(posedge \clk ) begin
        s80_val_n28 <= s79_val_n28;
    end
    always @(posedge \clk ) begin
        s80_val_n29 <= s79_val_n29;
    end
    always @(posedge \clk ) begin
        s80_val_n30 <= s79_val_n30;
    end
    always @(posedge \clk ) begin
        s80_val_n31 <= s79_val_n31;
    end
    always @(posedge \clk ) begin
        s80_val_n32 <= s79_val_n32;
    end
    always @(posedge \clk ) begin
        s80_val_n33 <= s79_val_n33;
    end
    always @(posedge \clk ) begin
        s80_val_n34 <= s79_val_n34;
    end
    always @(posedge \clk ) begin
        s80_val_n35 <= s79_val_n35;
    end
    always @(posedge \clk ) begin
        s80_val_n36 <= s79_val_n36;
    end
    always @(posedge \clk ) begin
        s80_val_n37 <= s79_val_n37;
    end
    always @(posedge \clk ) begin
        s80_val_n38 <= s79_val_n38;
    end
    always @(posedge \clk ) begin
        \s81_val  <= \s80_val ;
    end
    always @(posedge \clk ) begin
        s81_val_n1 <= s80_val_n1;
    end
    always @(posedge \clk ) begin
        s81_val_n2 <= s80_val_n2;
    end
    always @(posedge \clk ) begin
        s81_val_n3 <= s80_val_n3;
    end
    always @(posedge \clk ) begin
        s81_val_n4 <= s80_val_n4;
    end
    always @(posedge \clk ) begin
        s81_val_n5 <= s80_val_n5;
    end
    always @(posedge \clk ) begin
        s81_val_n6 <= s80_val_n6;
    end
    always @(posedge \clk ) begin
        s81_val_n7 <= s80_val_n7;
    end
    always @(posedge \clk ) begin
        s81_val_n8 <= s80_val_n8;
    end
    always @(posedge \clk ) begin
        s81_val_n9 <= s80_val_n9;
    end
    always @(posedge \clk ) begin
        s81_val_n10 <= s80_val_n10;
    end
    always @(posedge \clk ) begin
        s81_val_n11 <= s80_val_n11;
    end
    always @(posedge \clk ) begin
        s81_val_n12 <= s80_val_n12;
    end
    always @(posedge \clk ) begin
        s81_val_n13 <= s80_val_n13;
    end
    always @(posedge \clk ) begin
        s81_val_n14 <= s80_val_n14;
    end
    always @(posedge \clk ) begin
        s81_val_n15 <= s80_val_n15;
    end
    always @(posedge \clk ) begin
        s81_val_n16 <= s80_val_n16;
    end
    always @(posedge \clk ) begin
        s81_val_n17 <= s80_val_n17;
    end
    always @(posedge \clk ) begin
        s81_val_n18 <= s80_val_n18;
    end
    always @(posedge \clk ) begin
        s81_val_n19 <= s80_val_n19;
    end
    always @(posedge \clk ) begin
        s81_val_n20 <= s80_val_n20;
    end
    always @(posedge \clk ) begin
        s81_val_n21 <= s80_val_n21;
    end
    always @(posedge \clk ) begin
        s81_val_n22 <= s80_val_n22;
    end
    always @(posedge \clk ) begin
        s81_val_n23 <= s80_val_n23;
    end
    always @(posedge \clk ) begin
        s81_val_n24 <= s80_val_n24;
    end
    always @(posedge \clk ) begin
        s81_val_n25 <= s80_val_n25;
    end
    always @(posedge \clk ) begin
        s81_val_n26 <= s80_val_n26;
    end
    always @(posedge \clk ) begin
        s81_val_n27 <= s80_val_n27;
    end
    always @(posedge \clk ) begin
        s81_val_n28 <= s80_val_n28;
    end
    always @(posedge \clk ) begin
        s81_val_n29 <= s80_val_n29;
    end
    always @(posedge \clk ) begin
        s81_val_n30 <= s80_val_n30;
    end
    always @(posedge \clk ) begin
        s81_val_n31 <= s80_val_n31;
    end
    always @(posedge \clk ) begin
        s81_val_n32 <= s80_val_n32;
    end
    always @(posedge \clk ) begin
        s81_val_n33 <= s80_val_n33;
    end
    always @(posedge \clk ) begin
        s81_val_n34 <= s80_val_n34;
    end
    always @(posedge \clk ) begin
        s81_val_n35 <= s80_val_n35;
    end
    always @(posedge \clk ) begin
        s81_val_n36 <= s80_val_n36;
    end
    always @(posedge \clk ) begin
        s81_val_n37 <= s80_val_n37;
    end
    always @(posedge \clk ) begin
        s81_val_n38 <= s80_val_n38;
    end
    always @(posedge \clk ) begin
        s81_val_n39 <= val_n39;
    end
    always @(posedge \clk ) begin
        \s82_val  <= \s81_val ;
    end
    always @(posedge \clk ) begin
        s82_val_n1 <= s81_val_n1;
    end
    always @(posedge \clk ) begin
        s82_val_n2 <= s81_val_n2;
    end
    always @(posedge \clk ) begin
        s82_val_n3 <= s81_val_n3;
    end
    always @(posedge \clk ) begin
        s82_val_n4 <= s81_val_n4;
    end
    always @(posedge \clk ) begin
        s82_val_n5 <= s81_val_n5;
    end
    always @(posedge \clk ) begin
        s82_val_n6 <= s81_val_n6;
    end
    always @(posedge \clk ) begin
        s82_val_n7 <= s81_val_n7;
    end
    always @(posedge \clk ) begin
        s82_val_n8 <= s81_val_n8;
    end
    always @(posedge \clk ) begin
        s82_val_n9 <= s81_val_n9;
    end
    always @(posedge \clk ) begin
        s82_val_n10 <= s81_val_n10;
    end
    always @(posedge \clk ) begin
        s82_val_n11 <= s81_val_n11;
    end
    always @(posedge \clk ) begin
        s82_val_n12 <= s81_val_n12;
    end
    always @(posedge \clk ) begin
        s82_val_n13 <= s81_val_n13;
    end
    always @(posedge \clk ) begin
        s82_val_n14 <= s81_val_n14;
    end
    always @(posedge \clk ) begin
        s82_val_n15 <= s81_val_n15;
    end
    always @(posedge \clk ) begin
        s82_val_n16 <= s81_val_n16;
    end
    always @(posedge \clk ) begin
        s82_val_n17 <= s81_val_n17;
    end
    always @(posedge \clk ) begin
        s82_val_n18 <= s81_val_n18;
    end
    always @(posedge \clk ) begin
        s82_val_n19 <= s81_val_n19;
    end
    always @(posedge \clk ) begin
        s82_val_n20 <= s81_val_n20;
    end
    always @(posedge \clk ) begin
        s82_val_n21 <= s81_val_n21;
    end
    always @(posedge \clk ) begin
        s82_val_n22 <= s81_val_n22;
    end
    always @(posedge \clk ) begin
        s82_val_n23 <= s81_val_n23;
    end
    always @(posedge \clk ) begin
        s82_val_n24 <= s81_val_n24;
    end
    always @(posedge \clk ) begin
        s82_val_n25 <= s81_val_n25;
    end
    always @(posedge \clk ) begin
        s82_val_n26 <= s81_val_n26;
    end
    always @(posedge \clk ) begin
        s82_val_n27 <= s81_val_n27;
    end
    always @(posedge \clk ) begin
        s82_val_n28 <= s81_val_n28;
    end
    always @(posedge \clk ) begin
        s82_val_n29 <= s81_val_n29;
    end
    always @(posedge \clk ) begin
        s82_val_n30 <= s81_val_n30;
    end
    always @(posedge \clk ) begin
        s82_val_n31 <= s81_val_n31;
    end
    always @(posedge \clk ) begin
        s82_val_n32 <= s81_val_n32;
    end
    always @(posedge \clk ) begin
        s82_val_n33 <= s81_val_n33;
    end
    always @(posedge \clk ) begin
        s82_val_n34 <= s81_val_n34;
    end
    always @(posedge \clk ) begin
        s82_val_n35 <= s81_val_n35;
    end
    always @(posedge \clk ) begin
        s82_val_n36 <= s81_val_n36;
    end
    always @(posedge \clk ) begin
        s82_val_n37 <= s81_val_n37;
    end
    always @(posedge \clk ) begin
        s82_val_n38 <= s81_val_n38;
    end
    always @(posedge \clk ) begin
        s82_val_n39 <= s81_val_n39;
    end
    always @(posedge \clk ) begin
        \s83_val  <= \s82_val ;
    end
    always @(posedge \clk ) begin
        s83_val_n1 <= s82_val_n1;
    end
    always @(posedge \clk ) begin
        s83_val_n2 <= s82_val_n2;
    end
    always @(posedge \clk ) begin
        s83_val_n3 <= s82_val_n3;
    end
    always @(posedge \clk ) begin
        s83_val_n4 <= s82_val_n4;
    end
    always @(posedge \clk ) begin
        s83_val_n5 <= s82_val_n5;
    end
    always @(posedge \clk ) begin
        s83_val_n6 <= s82_val_n6;
    end
    always @(posedge \clk ) begin
        s83_val_n7 <= s82_val_n7;
    end
    always @(posedge \clk ) begin
        s83_val_n8 <= s82_val_n8;
    end
    always @(posedge \clk ) begin
        s83_val_n9 <= s82_val_n9;
    end
    always @(posedge \clk ) begin
        s83_val_n10 <= s82_val_n10;
    end
    always @(posedge \clk ) begin
        s83_val_n11 <= s82_val_n11;
    end
    always @(posedge \clk ) begin
        s83_val_n12 <= s82_val_n12;
    end
    always @(posedge \clk ) begin
        s83_val_n13 <= s82_val_n13;
    end
    always @(posedge \clk ) begin
        s83_val_n14 <= s82_val_n14;
    end
    always @(posedge \clk ) begin
        s83_val_n15 <= s82_val_n15;
    end
    always @(posedge \clk ) begin
        s83_val_n16 <= s82_val_n16;
    end
    always @(posedge \clk ) begin
        s83_val_n17 <= s82_val_n17;
    end
    always @(posedge \clk ) begin
        s83_val_n18 <= s82_val_n18;
    end
    always @(posedge \clk ) begin
        s83_val_n19 <= s82_val_n19;
    end
    always @(posedge \clk ) begin
        s83_val_n20 <= s82_val_n20;
    end
    always @(posedge \clk ) begin
        s83_val_n21 <= s82_val_n21;
    end
    always @(posedge \clk ) begin
        s83_val_n22 <= s82_val_n22;
    end
    always @(posedge \clk ) begin
        s83_val_n23 <= s82_val_n23;
    end
    always @(posedge \clk ) begin
        s83_val_n24 <= s82_val_n24;
    end
    always @(posedge \clk ) begin
        s83_val_n25 <= s82_val_n25;
    end
    always @(posedge \clk ) begin
        s83_val_n26 <= s82_val_n26;
    end
    always @(posedge \clk ) begin
        s83_val_n27 <= s82_val_n27;
    end
    always @(posedge \clk ) begin
        s83_val_n28 <= s82_val_n28;
    end
    always @(posedge \clk ) begin
        s83_val_n29 <= s82_val_n29;
    end
    always @(posedge \clk ) begin
        s83_val_n30 <= s82_val_n30;
    end
    always @(posedge \clk ) begin
        s83_val_n31 <= s82_val_n31;
    end
    always @(posedge \clk ) begin
        s83_val_n32 <= s82_val_n32;
    end
    always @(posedge \clk ) begin
        s83_val_n33 <= s82_val_n33;
    end
    always @(posedge \clk ) begin
        s83_val_n34 <= s82_val_n34;
    end
    always @(posedge \clk ) begin
        s83_val_n35 <= s82_val_n35;
    end
    always @(posedge \clk ) begin
        s83_val_n36 <= s82_val_n36;
    end
    always @(posedge \clk ) begin
        s83_val_n37 <= s82_val_n37;
    end
    always @(posedge \clk ) begin
        s83_val_n38 <= s82_val_n38;
    end
    always @(posedge \clk ) begin
        s83_val_n39 <= s82_val_n39;
    end
    always @(posedge \clk ) begin
        s83_val_n40 <= val_n40;
    end
    always @(posedge \clk ) begin
        \s84_val  <= \s83_val ;
    end
    always @(posedge \clk ) begin
        s84_val_n1 <= s83_val_n1;
    end
    always @(posedge \clk ) begin
        s84_val_n2 <= s83_val_n2;
    end
    always @(posedge \clk ) begin
        s84_val_n3 <= s83_val_n3;
    end
    always @(posedge \clk ) begin
        s84_val_n4 <= s83_val_n4;
    end
    always @(posedge \clk ) begin
        s84_val_n5 <= s83_val_n5;
    end
    always @(posedge \clk ) begin
        s84_val_n6 <= s83_val_n6;
    end
    always @(posedge \clk ) begin
        s84_val_n7 <= s83_val_n7;
    end
    always @(posedge \clk ) begin
        s84_val_n8 <= s83_val_n8;
    end
    always @(posedge \clk ) begin
        s84_val_n9 <= s83_val_n9;
    end
    always @(posedge \clk ) begin
        s84_val_n10 <= s83_val_n10;
    end
    always @(posedge \clk ) begin
        s84_val_n11 <= s83_val_n11;
    end
    always @(posedge \clk ) begin
        s84_val_n12 <= s83_val_n12;
    end
    always @(posedge \clk ) begin
        s84_val_n13 <= s83_val_n13;
    end
    always @(posedge \clk ) begin
        s84_val_n14 <= s83_val_n14;
    end
    always @(posedge \clk ) begin
        s84_val_n15 <= s83_val_n15;
    end
    always @(posedge \clk ) begin
        s84_val_n16 <= s83_val_n16;
    end
    always @(posedge \clk ) begin
        s84_val_n17 <= s83_val_n17;
    end
    always @(posedge \clk ) begin
        s84_val_n18 <= s83_val_n18;
    end
    always @(posedge \clk ) begin
        s84_val_n19 <= s83_val_n19;
    end
    always @(posedge \clk ) begin
        s84_val_n20 <= s83_val_n20;
    end
    always @(posedge \clk ) begin
        s84_val_n21 <= s83_val_n21;
    end
    always @(posedge \clk ) begin
        s84_val_n22 <= s83_val_n22;
    end
    always @(posedge \clk ) begin
        s84_val_n23 <= s83_val_n23;
    end
    always @(posedge \clk ) begin
        s84_val_n24 <= s83_val_n24;
    end
    always @(posedge \clk ) begin
        s84_val_n25 <= s83_val_n25;
    end
    always @(posedge \clk ) begin
        s84_val_n26 <= s83_val_n26;
    end
    always @(posedge \clk ) begin
        s84_val_n27 <= s83_val_n27;
    end
    always @(posedge \clk ) begin
        s84_val_n28 <= s83_val_n28;
    end
    always @(posedge \clk ) begin
        s84_val_n29 <= s83_val_n29;
    end
    always @(posedge \clk ) begin
        s84_val_n30 <= s83_val_n30;
    end
    always @(posedge \clk ) begin
        s84_val_n31 <= s83_val_n31;
    end
    always @(posedge \clk ) begin
        s84_val_n32 <= s83_val_n32;
    end
    always @(posedge \clk ) begin
        s84_val_n33 <= s83_val_n33;
    end
    always @(posedge \clk ) begin
        s84_val_n34 <= s83_val_n34;
    end
    always @(posedge \clk ) begin
        s84_val_n35 <= s83_val_n35;
    end
    always @(posedge \clk ) begin
        s84_val_n36 <= s83_val_n36;
    end
    always @(posedge \clk ) begin
        s84_val_n37 <= s83_val_n37;
    end
    always @(posedge \clk ) begin
        s84_val_n38 <= s83_val_n38;
    end
    always @(posedge \clk ) begin
        s84_val_n39 <= s83_val_n39;
    end
    always @(posedge \clk ) begin
        s84_val_n40 <= s83_val_n40;
    end
    always @(posedge \clk ) begin
        \s85_val  <= \s84_val ;
    end
    always @(posedge \clk ) begin
        s85_val_n1 <= s84_val_n1;
    end
    always @(posedge \clk ) begin
        s85_val_n2 <= s84_val_n2;
    end
    always @(posedge \clk ) begin
        s85_val_n3 <= s84_val_n3;
    end
    always @(posedge \clk ) begin
        s85_val_n4 <= s84_val_n4;
    end
    always @(posedge \clk ) begin
        s85_val_n5 <= s84_val_n5;
    end
    always @(posedge \clk ) begin
        s85_val_n6 <= s84_val_n6;
    end
    always @(posedge \clk ) begin
        s85_val_n7 <= s84_val_n7;
    end
    always @(posedge \clk ) begin
        s85_val_n8 <= s84_val_n8;
    end
    always @(posedge \clk ) begin
        s85_val_n9 <= s84_val_n9;
    end
    always @(posedge \clk ) begin
        s85_val_n10 <= s84_val_n10;
    end
    always @(posedge \clk ) begin
        s85_val_n11 <= s84_val_n11;
    end
    always @(posedge \clk ) begin
        s85_val_n12 <= s84_val_n12;
    end
    always @(posedge \clk ) begin
        s85_val_n13 <= s84_val_n13;
    end
    always @(posedge \clk ) begin
        s85_val_n14 <= s84_val_n14;
    end
    always @(posedge \clk ) begin
        s85_val_n15 <= s84_val_n15;
    end
    always @(posedge \clk ) begin
        s85_val_n16 <= s84_val_n16;
    end
    always @(posedge \clk ) begin
        s85_val_n17 <= s84_val_n17;
    end
    always @(posedge \clk ) begin
        s85_val_n18 <= s84_val_n18;
    end
    always @(posedge \clk ) begin
        s85_val_n19 <= s84_val_n19;
    end
    always @(posedge \clk ) begin
        s85_val_n20 <= s84_val_n20;
    end
    always @(posedge \clk ) begin
        s85_val_n21 <= s84_val_n21;
    end
    always @(posedge \clk ) begin
        s85_val_n22 <= s84_val_n22;
    end
    always @(posedge \clk ) begin
        s85_val_n23 <= s84_val_n23;
    end
    always @(posedge \clk ) begin
        s85_val_n24 <= s84_val_n24;
    end
    always @(posedge \clk ) begin
        s85_val_n25 <= s84_val_n25;
    end
    always @(posedge \clk ) begin
        s85_val_n26 <= s84_val_n26;
    end
    always @(posedge \clk ) begin
        s85_val_n27 <= s84_val_n27;
    end
    always @(posedge \clk ) begin
        s85_val_n28 <= s84_val_n28;
    end
    always @(posedge \clk ) begin
        s85_val_n29 <= s84_val_n29;
    end
    always @(posedge \clk ) begin
        s85_val_n30 <= s84_val_n30;
    end
    always @(posedge \clk ) begin
        s85_val_n31 <= s84_val_n31;
    end
    always @(posedge \clk ) begin
        s85_val_n32 <= s84_val_n32;
    end
    always @(posedge \clk ) begin
        s85_val_n33 <= s84_val_n33;
    end
    always @(posedge \clk ) begin
        s85_val_n34 <= s84_val_n34;
    end
    always @(posedge \clk ) begin
        s85_val_n35 <= s84_val_n35;
    end
    always @(posedge \clk ) begin
        s85_val_n36 <= s84_val_n36;
    end
    always @(posedge \clk ) begin
        s85_val_n37 <= s84_val_n37;
    end
    always @(posedge \clk ) begin
        s85_val_n38 <= s84_val_n38;
    end
    always @(posedge \clk ) begin
        s85_val_n39 <= s84_val_n39;
    end
    always @(posedge \clk ) begin
        s85_val_n40 <= s84_val_n40;
    end
    always @(posedge \clk ) begin
        s85_val_n41 <= val_n41;
    end
    always @(posedge \clk ) begin
        \s86_val  <= \s85_val ;
    end
    always @(posedge \clk ) begin
        s86_val_n1 <= s85_val_n1;
    end
    always @(posedge \clk ) begin
        s86_val_n2 <= s85_val_n2;
    end
    always @(posedge \clk ) begin
        s86_val_n3 <= s85_val_n3;
    end
    always @(posedge \clk ) begin
        s86_val_n4 <= s85_val_n4;
    end
    always @(posedge \clk ) begin
        s86_val_n5 <= s85_val_n5;
    end
    always @(posedge \clk ) begin
        s86_val_n6 <= s85_val_n6;
    end
    always @(posedge \clk ) begin
        s86_val_n7 <= s85_val_n7;
    end
    always @(posedge \clk ) begin
        s86_val_n8 <= s85_val_n8;
    end
    always @(posedge \clk ) begin
        s86_val_n9 <= s85_val_n9;
    end
    always @(posedge \clk ) begin
        s86_val_n10 <= s85_val_n10;
    end
    always @(posedge \clk ) begin
        s86_val_n11 <= s85_val_n11;
    end
    always @(posedge \clk ) begin
        s86_val_n12 <= s85_val_n12;
    end
    always @(posedge \clk ) begin
        s86_val_n13 <= s85_val_n13;
    end
    always @(posedge \clk ) begin
        s86_val_n14 <= s85_val_n14;
    end
    always @(posedge \clk ) begin
        s86_val_n15 <= s85_val_n15;
    end
    always @(posedge \clk ) begin
        s86_val_n16 <= s85_val_n16;
    end
    always @(posedge \clk ) begin
        s86_val_n17 <= s85_val_n17;
    end
    always @(posedge \clk ) begin
        s86_val_n18 <= s85_val_n18;
    end
    always @(posedge \clk ) begin
        s86_val_n19 <= s85_val_n19;
    end
    always @(posedge \clk ) begin
        s86_val_n20 <= s85_val_n20;
    end
    always @(posedge \clk ) begin
        s86_val_n21 <= s85_val_n21;
    end
    always @(posedge \clk ) begin
        s86_val_n22 <= s85_val_n22;
    end
    always @(posedge \clk ) begin
        s86_val_n23 <= s85_val_n23;
    end
    always @(posedge \clk ) begin
        s86_val_n24 <= s85_val_n24;
    end
    always @(posedge \clk ) begin
        s86_val_n25 <= s85_val_n25;
    end
    always @(posedge \clk ) begin
        s86_val_n26 <= s85_val_n26;
    end
    always @(posedge \clk ) begin
        s86_val_n27 <= s85_val_n27;
    end
    always @(posedge \clk ) begin
        s86_val_n28 <= s85_val_n28;
    end
    always @(posedge \clk ) begin
        s86_val_n29 <= s85_val_n29;
    end
    always @(posedge \clk ) begin
        s86_val_n30 <= s85_val_n30;
    end
    always @(posedge \clk ) begin
        s86_val_n31 <= s85_val_n31;
    end
    always @(posedge \clk ) begin
        s86_val_n32 <= s85_val_n32;
    end
    always @(posedge \clk ) begin
        s86_val_n33 <= s85_val_n33;
    end
    always @(posedge \clk ) begin
        s86_val_n34 <= s85_val_n34;
    end
    always @(posedge \clk ) begin
        s86_val_n35 <= s85_val_n35;
    end
    always @(posedge \clk ) begin
        s86_val_n36 <= s85_val_n36;
    end
    always @(posedge \clk ) begin
        s86_val_n37 <= s85_val_n37;
    end
    always @(posedge \clk ) begin
        s86_val_n38 <= s85_val_n38;
    end
    always @(posedge \clk ) begin
        s86_val_n39 <= s85_val_n39;
    end
    always @(posedge \clk ) begin
        s86_val_n40 <= s85_val_n40;
    end
    always @(posedge \clk ) begin
        s86_val_n41 <= s85_val_n41;
    end
    always @(posedge \clk ) begin
        \s87_val  <= \s86_val ;
    end
    always @(posedge \clk ) begin
        s87_val_n1 <= s86_val_n1;
    end
    always @(posedge \clk ) begin
        s87_val_n2 <= s86_val_n2;
    end
    always @(posedge \clk ) begin
        s87_val_n3 <= s86_val_n3;
    end
    always @(posedge \clk ) begin
        s87_val_n4 <= s86_val_n4;
    end
    always @(posedge \clk ) begin
        s87_val_n5 <= s86_val_n5;
    end
    always @(posedge \clk ) begin
        s87_val_n6 <= s86_val_n6;
    end
    always @(posedge \clk ) begin
        s87_val_n7 <= s86_val_n7;
    end
    always @(posedge \clk ) begin
        s87_val_n8 <= s86_val_n8;
    end
    always @(posedge \clk ) begin
        s87_val_n9 <= s86_val_n9;
    end
    always @(posedge \clk ) begin
        s87_val_n10 <= s86_val_n10;
    end
    always @(posedge \clk ) begin
        s87_val_n11 <= s86_val_n11;
    end
    always @(posedge \clk ) begin
        s87_val_n12 <= s86_val_n12;
    end
    always @(posedge \clk ) begin
        s87_val_n13 <= s86_val_n13;
    end
    always @(posedge \clk ) begin
        s87_val_n14 <= s86_val_n14;
    end
    always @(posedge \clk ) begin
        s87_val_n15 <= s86_val_n15;
    end
    always @(posedge \clk ) begin
        s87_val_n16 <= s86_val_n16;
    end
    always @(posedge \clk ) begin
        s87_val_n17 <= s86_val_n17;
    end
    always @(posedge \clk ) begin
        s87_val_n18 <= s86_val_n18;
    end
    always @(posedge \clk ) begin
        s87_val_n19 <= s86_val_n19;
    end
    always @(posedge \clk ) begin
        s87_val_n20 <= s86_val_n20;
    end
    always @(posedge \clk ) begin
        s87_val_n21 <= s86_val_n21;
    end
    always @(posedge \clk ) begin
        s87_val_n22 <= s86_val_n22;
    end
    always @(posedge \clk ) begin
        s87_val_n23 <= s86_val_n23;
    end
    always @(posedge \clk ) begin
        s87_val_n24 <= s86_val_n24;
    end
    always @(posedge \clk ) begin
        s87_val_n25 <= s86_val_n25;
    end
    always @(posedge \clk ) begin
        s87_val_n26 <= s86_val_n26;
    end
    always @(posedge \clk ) begin
        s87_val_n27 <= s86_val_n27;
    end
    always @(posedge \clk ) begin
        s87_val_n28 <= s86_val_n28;
    end
    always @(posedge \clk ) begin
        s87_val_n29 <= s86_val_n29;
    end
    always @(posedge \clk ) begin
        s87_val_n30 <= s86_val_n30;
    end
    always @(posedge \clk ) begin
        s87_val_n31 <= s86_val_n31;
    end
    always @(posedge \clk ) begin
        s87_val_n32 <= s86_val_n32;
    end
    always @(posedge \clk ) begin
        s87_val_n33 <= s86_val_n33;
    end
    always @(posedge \clk ) begin
        s87_val_n34 <= s86_val_n34;
    end
    always @(posedge \clk ) begin
        s87_val_n35 <= s86_val_n35;
    end
    always @(posedge \clk ) begin
        s87_val_n36 <= s86_val_n36;
    end
    always @(posedge \clk ) begin
        s87_val_n37 <= s86_val_n37;
    end
    always @(posedge \clk ) begin
        s87_val_n38 <= s86_val_n38;
    end
    always @(posedge \clk ) begin
        s87_val_n39 <= s86_val_n39;
    end
    always @(posedge \clk ) begin
        s87_val_n40 <= s86_val_n40;
    end
    always @(posedge \clk ) begin
        s87_val_n41 <= s86_val_n41;
    end
    always @(posedge \clk ) begin
        s87_val_n42 <= val_n42;
    end
    always @(posedge \clk ) begin
        \s88_val  <= \s87_val ;
    end
    always @(posedge \clk ) begin
        s88_val_n1 <= s87_val_n1;
    end
    always @(posedge \clk ) begin
        s88_val_n2 <= s87_val_n2;
    end
    always @(posedge \clk ) begin
        s88_val_n3 <= s87_val_n3;
    end
    always @(posedge \clk ) begin
        s88_val_n4 <= s87_val_n4;
    end
    always @(posedge \clk ) begin
        s88_val_n5 <= s87_val_n5;
    end
    always @(posedge \clk ) begin
        s88_val_n6 <= s87_val_n6;
    end
    always @(posedge \clk ) begin
        s88_val_n7 <= s87_val_n7;
    end
    always @(posedge \clk ) begin
        s88_val_n8 <= s87_val_n8;
    end
    always @(posedge \clk ) begin
        s88_val_n9 <= s87_val_n9;
    end
    always @(posedge \clk ) begin
        s88_val_n10 <= s87_val_n10;
    end
    always @(posedge \clk ) begin
        s88_val_n11 <= s87_val_n11;
    end
    always @(posedge \clk ) begin
        s88_val_n12 <= s87_val_n12;
    end
    always @(posedge \clk ) begin
        s88_val_n13 <= s87_val_n13;
    end
    always @(posedge \clk ) begin
        s88_val_n14 <= s87_val_n14;
    end
    always @(posedge \clk ) begin
        s88_val_n15 <= s87_val_n15;
    end
    always @(posedge \clk ) begin
        s88_val_n16 <= s87_val_n16;
    end
    always @(posedge \clk ) begin
        s88_val_n17 <= s87_val_n17;
    end
    always @(posedge \clk ) begin
        s88_val_n18 <= s87_val_n18;
    end
    always @(posedge \clk ) begin
        s88_val_n19 <= s87_val_n19;
    end
    always @(posedge \clk ) begin
        s88_val_n20 <= s87_val_n20;
    end
    always @(posedge \clk ) begin
        s88_val_n21 <= s87_val_n21;
    end
    always @(posedge \clk ) begin
        s88_val_n22 <= s87_val_n22;
    end
    always @(posedge \clk ) begin
        s88_val_n23 <= s87_val_n23;
    end
    always @(posedge \clk ) begin
        s88_val_n24 <= s87_val_n24;
    end
    always @(posedge \clk ) begin
        s88_val_n25 <= s87_val_n25;
    end
    always @(posedge \clk ) begin
        s88_val_n26 <= s87_val_n26;
    end
    always @(posedge \clk ) begin
        s88_val_n27 <= s87_val_n27;
    end
    always @(posedge \clk ) begin
        s88_val_n28 <= s87_val_n28;
    end
    always @(posedge \clk ) begin
        s88_val_n29 <= s87_val_n29;
    end
    always @(posedge \clk ) begin
        s88_val_n30 <= s87_val_n30;
    end
    always @(posedge \clk ) begin
        s88_val_n31 <= s87_val_n31;
    end
    always @(posedge \clk ) begin
        s88_val_n32 <= s87_val_n32;
    end
    always @(posedge \clk ) begin
        s88_val_n33 <= s87_val_n33;
    end
    always @(posedge \clk ) begin
        s88_val_n34 <= s87_val_n34;
    end
    always @(posedge \clk ) begin
        s88_val_n35 <= s87_val_n35;
    end
    always @(posedge \clk ) begin
        s88_val_n36 <= s87_val_n36;
    end
    always @(posedge \clk ) begin
        s88_val_n37 <= s87_val_n37;
    end
    always @(posedge \clk ) begin
        s88_val_n38 <= s87_val_n38;
    end
    always @(posedge \clk ) begin
        s88_val_n39 <= s87_val_n39;
    end
    always @(posedge \clk ) begin
        s88_val_n40 <= s87_val_n40;
    end
    always @(posedge \clk ) begin
        s88_val_n41 <= s87_val_n41;
    end
    always @(posedge \clk ) begin
        s88_val_n42 <= s87_val_n42;
    end
    always @(posedge \clk ) begin
        \s89_val  <= \s88_val ;
    end
    always @(posedge \clk ) begin
        s89_val_n1 <= s88_val_n1;
    end
    always @(posedge \clk ) begin
        s89_val_n2 <= s88_val_n2;
    end
    always @(posedge \clk ) begin
        s89_val_n3 <= s88_val_n3;
    end
    always @(posedge \clk ) begin
        s89_val_n4 <= s88_val_n4;
    end
    always @(posedge \clk ) begin
        s89_val_n5 <= s88_val_n5;
    end
    always @(posedge \clk ) begin
        s89_val_n6 <= s88_val_n6;
    end
    always @(posedge \clk ) begin
        s89_val_n7 <= s88_val_n7;
    end
    always @(posedge \clk ) begin
        s89_val_n8 <= s88_val_n8;
    end
    always @(posedge \clk ) begin
        s89_val_n9 <= s88_val_n9;
    end
    always @(posedge \clk ) begin
        s89_val_n10 <= s88_val_n10;
    end
    always @(posedge \clk ) begin
        s89_val_n11 <= s88_val_n11;
    end
    always @(posedge \clk ) begin
        s89_val_n12 <= s88_val_n12;
    end
    always @(posedge \clk ) begin
        s89_val_n13 <= s88_val_n13;
    end
    always @(posedge \clk ) begin
        s89_val_n14 <= s88_val_n14;
    end
    always @(posedge \clk ) begin
        s89_val_n15 <= s88_val_n15;
    end
    always @(posedge \clk ) begin
        s89_val_n16 <= s88_val_n16;
    end
    always @(posedge \clk ) begin
        s89_val_n17 <= s88_val_n17;
    end
    always @(posedge \clk ) begin
        s89_val_n18 <= s88_val_n18;
    end
    always @(posedge \clk ) begin
        s89_val_n19 <= s88_val_n19;
    end
    always @(posedge \clk ) begin
        s89_val_n20 <= s88_val_n20;
    end
    always @(posedge \clk ) begin
        s89_val_n21 <= s88_val_n21;
    end
    always @(posedge \clk ) begin
        s89_val_n22 <= s88_val_n22;
    end
    always @(posedge \clk ) begin
        s89_val_n23 <= s88_val_n23;
    end
    always @(posedge \clk ) begin
        s89_val_n24 <= s88_val_n24;
    end
    always @(posedge \clk ) begin
        s89_val_n25 <= s88_val_n25;
    end
    always @(posedge \clk ) begin
        s89_val_n26 <= s88_val_n26;
    end
    always @(posedge \clk ) begin
        s89_val_n27 <= s88_val_n27;
    end
    always @(posedge \clk ) begin
        s89_val_n28 <= s88_val_n28;
    end
    always @(posedge \clk ) begin
        s89_val_n29 <= s88_val_n29;
    end
    always @(posedge \clk ) begin
        s89_val_n30 <= s88_val_n30;
    end
    always @(posedge \clk ) begin
        s89_val_n31 <= s88_val_n31;
    end
    always @(posedge \clk ) begin
        s89_val_n32 <= s88_val_n32;
    end
    always @(posedge \clk ) begin
        s89_val_n33 <= s88_val_n33;
    end
    always @(posedge \clk ) begin
        s89_val_n34 <= s88_val_n34;
    end
    always @(posedge \clk ) begin
        s89_val_n35 <= s88_val_n35;
    end
    always @(posedge \clk ) begin
        s89_val_n36 <= s88_val_n36;
    end
    always @(posedge \clk ) begin
        s89_val_n37 <= s88_val_n37;
    end
    always @(posedge \clk ) begin
        s89_val_n38 <= s88_val_n38;
    end
    always @(posedge \clk ) begin
        s89_val_n39 <= s88_val_n39;
    end
    always @(posedge \clk ) begin
        s89_val_n40 <= s88_val_n40;
    end
    always @(posedge \clk ) begin
        s89_val_n41 <= s88_val_n41;
    end
    always @(posedge \clk ) begin
        s89_val_n42 <= s88_val_n42;
    end
    always @(posedge \clk ) begin
        s89_val_n43 <= val_n43;
    end
    always @(posedge \clk ) begin
        \s90_val  <= \s89_val ;
    end
    always @(posedge \clk ) begin
        s90_val_n1 <= s89_val_n1;
    end
    always @(posedge \clk ) begin
        s90_val_n2 <= s89_val_n2;
    end
    always @(posedge \clk ) begin
        s90_val_n3 <= s89_val_n3;
    end
    always @(posedge \clk ) begin
        s90_val_n4 <= s89_val_n4;
    end
    always @(posedge \clk ) begin
        s90_val_n5 <= s89_val_n5;
    end
    always @(posedge \clk ) begin
        s90_val_n6 <= s89_val_n6;
    end
    always @(posedge \clk ) begin
        s90_val_n7 <= s89_val_n7;
    end
    always @(posedge \clk ) begin
        s90_val_n8 <= s89_val_n8;
    end
    always @(posedge \clk ) begin
        s90_val_n9 <= s89_val_n9;
    end
    always @(posedge \clk ) begin
        s90_val_n10 <= s89_val_n10;
    end
    always @(posedge \clk ) begin
        s90_val_n11 <= s89_val_n11;
    end
    always @(posedge \clk ) begin
        s90_val_n12 <= s89_val_n12;
    end
    always @(posedge \clk ) begin
        s90_val_n13 <= s89_val_n13;
    end
    always @(posedge \clk ) begin
        s90_val_n14 <= s89_val_n14;
    end
    always @(posedge \clk ) begin
        s90_val_n15 <= s89_val_n15;
    end
    always @(posedge \clk ) begin
        s90_val_n16 <= s89_val_n16;
    end
    always @(posedge \clk ) begin
        s90_val_n17 <= s89_val_n17;
    end
    always @(posedge \clk ) begin
        s90_val_n18 <= s89_val_n18;
    end
    always @(posedge \clk ) begin
        s90_val_n19 <= s89_val_n19;
    end
    always @(posedge \clk ) begin
        s90_val_n20 <= s89_val_n20;
    end
    always @(posedge \clk ) begin
        s90_val_n21 <= s89_val_n21;
    end
    always @(posedge \clk ) begin
        s90_val_n22 <= s89_val_n22;
    end
    always @(posedge \clk ) begin
        s90_val_n23 <= s89_val_n23;
    end
    always @(posedge \clk ) begin
        s90_val_n24 <= s89_val_n24;
    end
    always @(posedge \clk ) begin
        s90_val_n25 <= s89_val_n25;
    end
    always @(posedge \clk ) begin
        s90_val_n26 <= s89_val_n26;
    end
    always @(posedge \clk ) begin
        s90_val_n27 <= s89_val_n27;
    end
    always @(posedge \clk ) begin
        s90_val_n28 <= s89_val_n28;
    end
    always @(posedge \clk ) begin
        s90_val_n29 <= s89_val_n29;
    end
    always @(posedge \clk ) begin
        s90_val_n30 <= s89_val_n30;
    end
    always @(posedge \clk ) begin
        s90_val_n31 <= s89_val_n31;
    end
    always @(posedge \clk ) begin
        s90_val_n32 <= s89_val_n32;
    end
    always @(posedge \clk ) begin
        s90_val_n33 <= s89_val_n33;
    end
    always @(posedge \clk ) begin
        s90_val_n34 <= s89_val_n34;
    end
    always @(posedge \clk ) begin
        s90_val_n35 <= s89_val_n35;
    end
    always @(posedge \clk ) begin
        s90_val_n36 <= s89_val_n36;
    end
    always @(posedge \clk ) begin
        s90_val_n37 <= s89_val_n37;
    end
    always @(posedge \clk ) begin
        s90_val_n38 <= s89_val_n38;
    end
    always @(posedge \clk ) begin
        s90_val_n39 <= s89_val_n39;
    end
    always @(posedge \clk ) begin
        s90_val_n40 <= s89_val_n40;
    end
    always @(posedge \clk ) begin
        s90_val_n41 <= s89_val_n41;
    end
    always @(posedge \clk ) begin
        s90_val_n42 <= s89_val_n42;
    end
    always @(posedge \clk ) begin
        s90_val_n43 <= s89_val_n43;
    end
    always @(posedge \clk ) begin
        \s91_val  <= \s90_val ;
    end
    always @(posedge \clk ) begin
        s91_val_n1 <= s90_val_n1;
    end
    always @(posedge \clk ) begin
        s91_val_n2 <= s90_val_n2;
    end
    always @(posedge \clk ) begin
        s91_val_n3 <= s90_val_n3;
    end
    always @(posedge \clk ) begin
        s91_val_n4 <= s90_val_n4;
    end
    always @(posedge \clk ) begin
        s91_val_n5 <= s90_val_n5;
    end
    always @(posedge \clk ) begin
        s91_val_n6 <= s90_val_n6;
    end
    always @(posedge \clk ) begin
        s91_val_n7 <= s90_val_n7;
    end
    always @(posedge \clk ) begin
        s91_val_n8 <= s90_val_n8;
    end
    always @(posedge \clk ) begin
        s91_val_n9 <= s90_val_n9;
    end
    always @(posedge \clk ) begin
        s91_val_n10 <= s90_val_n10;
    end
    always @(posedge \clk ) begin
        s91_val_n11 <= s90_val_n11;
    end
    always @(posedge \clk ) begin
        s91_val_n12 <= s90_val_n12;
    end
    always @(posedge \clk ) begin
        s91_val_n13 <= s90_val_n13;
    end
    always @(posedge \clk ) begin
        s91_val_n14 <= s90_val_n14;
    end
    always @(posedge \clk ) begin
        s91_val_n15 <= s90_val_n15;
    end
    always @(posedge \clk ) begin
        s91_val_n16 <= s90_val_n16;
    end
    always @(posedge \clk ) begin
        s91_val_n17 <= s90_val_n17;
    end
    always @(posedge \clk ) begin
        s91_val_n18 <= s90_val_n18;
    end
    always @(posedge \clk ) begin
        s91_val_n19 <= s90_val_n19;
    end
    always @(posedge \clk ) begin
        s91_val_n20 <= s90_val_n20;
    end
    always @(posedge \clk ) begin
        s91_val_n21 <= s90_val_n21;
    end
    always @(posedge \clk ) begin
        s91_val_n22 <= s90_val_n22;
    end
    always @(posedge \clk ) begin
        s91_val_n23 <= s90_val_n23;
    end
    always @(posedge \clk ) begin
        s91_val_n24 <= s90_val_n24;
    end
    always @(posedge \clk ) begin
        s91_val_n25 <= s90_val_n25;
    end
    always @(posedge \clk ) begin
        s91_val_n26 <= s90_val_n26;
    end
    always @(posedge \clk ) begin
        s91_val_n27 <= s90_val_n27;
    end
    always @(posedge \clk ) begin
        s91_val_n28 <= s90_val_n28;
    end
    always @(posedge \clk ) begin
        s91_val_n29 <= s90_val_n29;
    end
    always @(posedge \clk ) begin
        s91_val_n30 <= s90_val_n30;
    end
    always @(posedge \clk ) begin
        s91_val_n31 <= s90_val_n31;
    end
    always @(posedge \clk ) begin
        s91_val_n32 <= s90_val_n32;
    end
    always @(posedge \clk ) begin
        s91_val_n33 <= s90_val_n33;
    end
    always @(posedge \clk ) begin
        s91_val_n34 <= s90_val_n34;
    end
    always @(posedge \clk ) begin
        s91_val_n35 <= s90_val_n35;
    end
    always @(posedge \clk ) begin
        s91_val_n36 <= s90_val_n36;
    end
    always @(posedge \clk ) begin
        s91_val_n37 <= s90_val_n37;
    end
    always @(posedge \clk ) begin
        s91_val_n38 <= s90_val_n38;
    end
    always @(posedge \clk ) begin
        s91_val_n39 <= s90_val_n39;
    end
    always @(posedge \clk ) begin
        s91_val_n40 <= s90_val_n40;
    end
    always @(posedge \clk ) begin
        s91_val_n41 <= s90_val_n41;
    end
    always @(posedge \clk ) begin
        s91_val_n42 <= s90_val_n42;
    end
    always @(posedge \clk ) begin
        s91_val_n43 <= s90_val_n43;
    end
    always @(posedge \clk ) begin
        s91_val_n44 <= val_n44;
    end
    always @(posedge \clk ) begin
        \s92_val  <= \s91_val ;
    end
    always @(posedge \clk ) begin
        s92_val_n1 <= s91_val_n1;
    end
    always @(posedge \clk ) begin
        s92_val_n2 <= s91_val_n2;
    end
    always @(posedge \clk ) begin
        s92_val_n3 <= s91_val_n3;
    end
    always @(posedge \clk ) begin
        s92_val_n4 <= s91_val_n4;
    end
    always @(posedge \clk ) begin
        s92_val_n5 <= s91_val_n5;
    end
    always @(posedge \clk ) begin
        s92_val_n6 <= s91_val_n6;
    end
    always @(posedge \clk ) begin
        s92_val_n7 <= s91_val_n7;
    end
    always @(posedge \clk ) begin
        s92_val_n8 <= s91_val_n8;
    end
    always @(posedge \clk ) begin
        s92_val_n9 <= s91_val_n9;
    end
    always @(posedge \clk ) begin
        s92_val_n10 <= s91_val_n10;
    end
    always @(posedge \clk ) begin
        s92_val_n11 <= s91_val_n11;
    end
    always @(posedge \clk ) begin
        s92_val_n12 <= s91_val_n12;
    end
    always @(posedge \clk ) begin
        s92_val_n13 <= s91_val_n13;
    end
    always @(posedge \clk ) begin
        s92_val_n14 <= s91_val_n14;
    end
    always @(posedge \clk ) begin
        s92_val_n15 <= s91_val_n15;
    end
    always @(posedge \clk ) begin
        s92_val_n16 <= s91_val_n16;
    end
    always @(posedge \clk ) begin
        s92_val_n17 <= s91_val_n17;
    end
    always @(posedge \clk ) begin
        s92_val_n18 <= s91_val_n18;
    end
    always @(posedge \clk ) begin
        s92_val_n19 <= s91_val_n19;
    end
    always @(posedge \clk ) begin
        s92_val_n20 <= s91_val_n20;
    end
    always @(posedge \clk ) begin
        s92_val_n21 <= s91_val_n21;
    end
    always @(posedge \clk ) begin
        s92_val_n22 <= s91_val_n22;
    end
    always @(posedge \clk ) begin
        s92_val_n23 <= s91_val_n23;
    end
    always @(posedge \clk ) begin
        s92_val_n24 <= s91_val_n24;
    end
    always @(posedge \clk ) begin
        s92_val_n25 <= s91_val_n25;
    end
    always @(posedge \clk ) begin
        s92_val_n26 <= s91_val_n26;
    end
    always @(posedge \clk ) begin
        s92_val_n27 <= s91_val_n27;
    end
    always @(posedge \clk ) begin
        s92_val_n28 <= s91_val_n28;
    end
    always @(posedge \clk ) begin
        s92_val_n29 <= s91_val_n29;
    end
    always @(posedge \clk ) begin
        s92_val_n30 <= s91_val_n30;
    end
    always @(posedge \clk ) begin
        s92_val_n31 <= s91_val_n31;
    end
    always @(posedge \clk ) begin
        s92_val_n32 <= s91_val_n32;
    end
    always @(posedge \clk ) begin
        s92_val_n33 <= s91_val_n33;
    end
    always @(posedge \clk ) begin
        s92_val_n34 <= s91_val_n34;
    end
    always @(posedge \clk ) begin
        s92_val_n35 <= s91_val_n35;
    end
    always @(posedge \clk ) begin
        s92_val_n36 <= s91_val_n36;
    end
    always @(posedge \clk ) begin
        s92_val_n37 <= s91_val_n37;
    end
    always @(posedge \clk ) begin
        s92_val_n38 <= s91_val_n38;
    end
    always @(posedge \clk ) begin
        s92_val_n39 <= s91_val_n39;
    end
    always @(posedge \clk ) begin
        s92_val_n40 <= s91_val_n40;
    end
    always @(posedge \clk ) begin
        s92_val_n41 <= s91_val_n41;
    end
    always @(posedge \clk ) begin
        s92_val_n42 <= s91_val_n42;
    end
    always @(posedge \clk ) begin
        s92_val_n43 <= s91_val_n43;
    end
    always @(posedge \clk ) begin
        s92_val_n44 <= s91_val_n44;
    end
    always @(posedge \clk ) begin
        \s93_val  <= \s92_val ;
    end
    always @(posedge \clk ) begin
        s93_val_n1 <= s92_val_n1;
    end
    always @(posedge \clk ) begin
        s93_val_n2 <= s92_val_n2;
    end
    always @(posedge \clk ) begin
        s93_val_n3 <= s92_val_n3;
    end
    always @(posedge \clk ) begin
        s93_val_n4 <= s92_val_n4;
    end
    always @(posedge \clk ) begin
        s93_val_n5 <= s92_val_n5;
    end
    always @(posedge \clk ) begin
        s93_val_n6 <= s92_val_n6;
    end
    always @(posedge \clk ) begin
        s93_val_n7 <= s92_val_n7;
    end
    always @(posedge \clk ) begin
        s93_val_n8 <= s92_val_n8;
    end
    always @(posedge \clk ) begin
        s93_val_n9 <= s92_val_n9;
    end
    always @(posedge \clk ) begin
        s93_val_n10 <= s92_val_n10;
    end
    always @(posedge \clk ) begin
        s93_val_n11 <= s92_val_n11;
    end
    always @(posedge \clk ) begin
        s93_val_n12 <= s92_val_n12;
    end
    always @(posedge \clk ) begin
        s93_val_n13 <= s92_val_n13;
    end
    always @(posedge \clk ) begin
        s93_val_n14 <= s92_val_n14;
    end
    always @(posedge \clk ) begin
        s93_val_n15 <= s92_val_n15;
    end
    always @(posedge \clk ) begin
        s93_val_n16 <= s92_val_n16;
    end
    always @(posedge \clk ) begin
        s93_val_n17 <= s92_val_n17;
    end
    always @(posedge \clk ) begin
        s93_val_n18 <= s92_val_n18;
    end
    always @(posedge \clk ) begin
        s93_val_n19 <= s92_val_n19;
    end
    always @(posedge \clk ) begin
        s93_val_n20 <= s92_val_n20;
    end
    always @(posedge \clk ) begin
        s93_val_n21 <= s92_val_n21;
    end
    always @(posedge \clk ) begin
        s93_val_n22 <= s92_val_n22;
    end
    always @(posedge \clk ) begin
        s93_val_n23 <= s92_val_n23;
    end
    always @(posedge \clk ) begin
        s93_val_n24 <= s92_val_n24;
    end
    always @(posedge \clk ) begin
        s93_val_n25 <= s92_val_n25;
    end
    always @(posedge \clk ) begin
        s93_val_n26 <= s92_val_n26;
    end
    always @(posedge \clk ) begin
        s93_val_n27 <= s92_val_n27;
    end
    always @(posedge \clk ) begin
        s93_val_n28 <= s92_val_n28;
    end
    always @(posedge \clk ) begin
        s93_val_n29 <= s92_val_n29;
    end
    always @(posedge \clk ) begin
        s93_val_n30 <= s92_val_n30;
    end
    always @(posedge \clk ) begin
        s93_val_n31 <= s92_val_n31;
    end
    always @(posedge \clk ) begin
        s93_val_n32 <= s92_val_n32;
    end
    always @(posedge \clk ) begin
        s93_val_n33 <= s92_val_n33;
    end
    always @(posedge \clk ) begin
        s93_val_n34 <= s92_val_n34;
    end
    always @(posedge \clk ) begin
        s93_val_n35 <= s92_val_n35;
    end
    always @(posedge \clk ) begin
        s93_val_n36 <= s92_val_n36;
    end
    always @(posedge \clk ) begin
        s93_val_n37 <= s92_val_n37;
    end
    always @(posedge \clk ) begin
        s93_val_n38 <= s92_val_n38;
    end
    always @(posedge \clk ) begin
        s93_val_n39 <= s92_val_n39;
    end
    always @(posedge \clk ) begin
        s93_val_n40 <= s92_val_n40;
    end
    always @(posedge \clk ) begin
        s93_val_n41 <= s92_val_n41;
    end
    always @(posedge \clk ) begin
        s93_val_n42 <= s92_val_n42;
    end
    always @(posedge \clk ) begin
        s93_val_n43 <= s92_val_n43;
    end
    always @(posedge \clk ) begin
        s93_val_n44 <= s92_val_n44;
    end
    always @(posedge \clk ) begin
        s93_val_n45 <= val_n45;
    end
    always @(posedge \clk ) begin
        \s94_val  <= \s93_val ;
    end
    always @(posedge \clk ) begin
        s94_val_n1 <= s93_val_n1;
    end
    always @(posedge \clk ) begin
        s94_val_n2 <= s93_val_n2;
    end
    always @(posedge \clk ) begin
        s94_val_n3 <= s93_val_n3;
    end
    always @(posedge \clk ) begin
        s94_val_n4 <= s93_val_n4;
    end
    always @(posedge \clk ) begin
        s94_val_n5 <= s93_val_n5;
    end
    always @(posedge \clk ) begin
        s94_val_n6 <= s93_val_n6;
    end
    always @(posedge \clk ) begin
        s94_val_n7 <= s93_val_n7;
    end
    always @(posedge \clk ) begin
        s94_val_n8 <= s93_val_n8;
    end
    always @(posedge \clk ) begin
        s94_val_n9 <= s93_val_n9;
    end
    always @(posedge \clk ) begin
        s94_val_n10 <= s93_val_n10;
    end
    always @(posedge \clk ) begin
        s94_val_n11 <= s93_val_n11;
    end
    always @(posedge \clk ) begin
        s94_val_n12 <= s93_val_n12;
    end
    always @(posedge \clk ) begin
        s94_val_n13 <= s93_val_n13;
    end
    always @(posedge \clk ) begin
        s94_val_n14 <= s93_val_n14;
    end
    always @(posedge \clk ) begin
        s94_val_n15 <= s93_val_n15;
    end
    always @(posedge \clk ) begin
        s94_val_n16 <= s93_val_n16;
    end
    always @(posedge \clk ) begin
        s94_val_n17 <= s93_val_n17;
    end
    always @(posedge \clk ) begin
        s94_val_n18 <= s93_val_n18;
    end
    always @(posedge \clk ) begin
        s94_val_n19 <= s93_val_n19;
    end
    always @(posedge \clk ) begin
        s94_val_n20 <= s93_val_n20;
    end
    always @(posedge \clk ) begin
        s94_val_n21 <= s93_val_n21;
    end
    always @(posedge \clk ) begin
        s94_val_n22 <= s93_val_n22;
    end
    always @(posedge \clk ) begin
        s94_val_n23 <= s93_val_n23;
    end
    always @(posedge \clk ) begin
        s94_val_n24 <= s93_val_n24;
    end
    always @(posedge \clk ) begin
        s94_val_n25 <= s93_val_n25;
    end
    always @(posedge \clk ) begin
        s94_val_n26 <= s93_val_n26;
    end
    always @(posedge \clk ) begin
        s94_val_n27 <= s93_val_n27;
    end
    always @(posedge \clk ) begin
        s94_val_n28 <= s93_val_n28;
    end
    always @(posedge \clk ) begin
        s94_val_n29 <= s93_val_n29;
    end
    always @(posedge \clk ) begin
        s94_val_n30 <= s93_val_n30;
    end
    always @(posedge \clk ) begin
        s94_val_n31 <= s93_val_n31;
    end
    always @(posedge \clk ) begin
        s94_val_n32 <= s93_val_n32;
    end
    always @(posedge \clk ) begin
        s94_val_n33 <= s93_val_n33;
    end
    always @(posedge \clk ) begin
        s94_val_n34 <= s93_val_n34;
    end
    always @(posedge \clk ) begin
        s94_val_n35 <= s93_val_n35;
    end
    always @(posedge \clk ) begin
        s94_val_n36 <= s93_val_n36;
    end
    always @(posedge \clk ) begin
        s94_val_n37 <= s93_val_n37;
    end
    always @(posedge \clk ) begin
        s94_val_n38 <= s93_val_n38;
    end
    always @(posedge \clk ) begin
        s94_val_n39 <= s93_val_n39;
    end
    always @(posedge \clk ) begin
        s94_val_n40 <= s93_val_n40;
    end
    always @(posedge \clk ) begin
        s94_val_n41 <= s93_val_n41;
    end
    always @(posedge \clk ) begin
        s94_val_n42 <= s93_val_n42;
    end
    always @(posedge \clk ) begin
        s94_val_n43 <= s93_val_n43;
    end
    always @(posedge \clk ) begin
        s94_val_n44 <= s93_val_n44;
    end
    always @(posedge \clk ) begin
        s94_val_n45 <= s93_val_n45;
    end
    always @(posedge \clk ) begin
        \s95_val  <= \s94_val ;
    end
    always @(posedge \clk ) begin
        s95_val_n1 <= s94_val_n1;
    end
    always @(posedge \clk ) begin
        s95_val_n2 <= s94_val_n2;
    end
    always @(posedge \clk ) begin
        s95_val_n3 <= s94_val_n3;
    end
    always @(posedge \clk ) begin
        s95_val_n4 <= s94_val_n4;
    end
    always @(posedge \clk ) begin
        s95_val_n5 <= s94_val_n5;
    end
    always @(posedge \clk ) begin
        s95_val_n6 <= s94_val_n6;
    end
    always @(posedge \clk ) begin
        s95_val_n7 <= s94_val_n7;
    end
    always @(posedge \clk ) begin
        s95_val_n8 <= s94_val_n8;
    end
    always @(posedge \clk ) begin
        s95_val_n9 <= s94_val_n9;
    end
    always @(posedge \clk ) begin
        s95_val_n10 <= s94_val_n10;
    end
    always @(posedge \clk ) begin
        s95_val_n11 <= s94_val_n11;
    end
    always @(posedge \clk ) begin
        s95_val_n12 <= s94_val_n12;
    end
    always @(posedge \clk ) begin
        s95_val_n13 <= s94_val_n13;
    end
    always @(posedge \clk ) begin
        s95_val_n14 <= s94_val_n14;
    end
    always @(posedge \clk ) begin
        s95_val_n15 <= s94_val_n15;
    end
    always @(posedge \clk ) begin
        s95_val_n16 <= s94_val_n16;
    end
    always @(posedge \clk ) begin
        s95_val_n17 <= s94_val_n17;
    end
    always @(posedge \clk ) begin
        s95_val_n18 <= s94_val_n18;
    end
    always @(posedge \clk ) begin
        s95_val_n19 <= s94_val_n19;
    end
    always @(posedge \clk ) begin
        s95_val_n20 <= s94_val_n20;
    end
    always @(posedge \clk ) begin
        s95_val_n21 <= s94_val_n21;
    end
    always @(posedge \clk ) begin
        s95_val_n22 <= s94_val_n22;
    end
    always @(posedge \clk ) begin
        s95_val_n23 <= s94_val_n23;
    end
    always @(posedge \clk ) begin
        s95_val_n24 <= s94_val_n24;
    end
    always @(posedge \clk ) begin
        s95_val_n25 <= s94_val_n25;
    end
    always @(posedge \clk ) begin
        s95_val_n26 <= s94_val_n26;
    end
    always @(posedge \clk ) begin
        s95_val_n27 <= s94_val_n27;
    end
    always @(posedge \clk ) begin
        s95_val_n28 <= s94_val_n28;
    end
    always @(posedge \clk ) begin
        s95_val_n29 <= s94_val_n29;
    end
    always @(posedge \clk ) begin
        s95_val_n30 <= s94_val_n30;
    end
    always @(posedge \clk ) begin
        s95_val_n31 <= s94_val_n31;
    end
    always @(posedge \clk ) begin
        s95_val_n32 <= s94_val_n32;
    end
    always @(posedge \clk ) begin
        s95_val_n33 <= s94_val_n33;
    end
    always @(posedge \clk ) begin
        s95_val_n34 <= s94_val_n34;
    end
    always @(posedge \clk ) begin
        s95_val_n35 <= s94_val_n35;
    end
    always @(posedge \clk ) begin
        s95_val_n36 <= s94_val_n36;
    end
    always @(posedge \clk ) begin
        s95_val_n37 <= s94_val_n37;
    end
    always @(posedge \clk ) begin
        s95_val_n38 <= s94_val_n38;
    end
    always @(posedge \clk ) begin
        s95_val_n39 <= s94_val_n39;
    end
    always @(posedge \clk ) begin
        s95_val_n40 <= s94_val_n40;
    end
    always @(posedge \clk ) begin
        s95_val_n41 <= s94_val_n41;
    end
    always @(posedge \clk ) begin
        s95_val_n42 <= s94_val_n42;
    end
    always @(posedge \clk ) begin
        s95_val_n43 <= s94_val_n43;
    end
    always @(posedge \clk ) begin
        s95_val_n44 <= s94_val_n44;
    end
    always @(posedge \clk ) begin
        s95_val_n45 <= s94_val_n45;
    end
    always @(posedge \clk ) begin
        s95_val_n46 <= val_n46;
    end
    always @(posedge \clk ) begin
        \s96_val  <= \s95_val ;
    end
    always @(posedge \clk ) begin
        s96_val_n1 <= s95_val_n1;
    end
    always @(posedge \clk ) begin
        s96_val_n2 <= s95_val_n2;
    end
    always @(posedge \clk ) begin
        s96_val_n3 <= s95_val_n3;
    end
    always @(posedge \clk ) begin
        s96_val_n4 <= s95_val_n4;
    end
    always @(posedge \clk ) begin
        s96_val_n5 <= s95_val_n5;
    end
    always @(posedge \clk ) begin
        s96_val_n6 <= s95_val_n6;
    end
    always @(posedge \clk ) begin
        s96_val_n7 <= s95_val_n7;
    end
    always @(posedge \clk ) begin
        s96_val_n8 <= s95_val_n8;
    end
    always @(posedge \clk ) begin
        s96_val_n9 <= s95_val_n9;
    end
    always @(posedge \clk ) begin
        s96_val_n10 <= s95_val_n10;
    end
    always @(posedge \clk ) begin
        s96_val_n11 <= s95_val_n11;
    end
    always @(posedge \clk ) begin
        s96_val_n12 <= s95_val_n12;
    end
    always @(posedge \clk ) begin
        s96_val_n13 <= s95_val_n13;
    end
    always @(posedge \clk ) begin
        s96_val_n14 <= s95_val_n14;
    end
    always @(posedge \clk ) begin
        s96_val_n15 <= s95_val_n15;
    end
    always @(posedge \clk ) begin
        s96_val_n16 <= s95_val_n16;
    end
    always @(posedge \clk ) begin
        s96_val_n17 <= s95_val_n17;
    end
    always @(posedge \clk ) begin
        s96_val_n18 <= s95_val_n18;
    end
    always @(posedge \clk ) begin
        s96_val_n19 <= s95_val_n19;
    end
    always @(posedge \clk ) begin
        s96_val_n20 <= s95_val_n20;
    end
    always @(posedge \clk ) begin
        s96_val_n21 <= s95_val_n21;
    end
    always @(posedge \clk ) begin
        s96_val_n22 <= s95_val_n22;
    end
    always @(posedge \clk ) begin
        s96_val_n23 <= s95_val_n23;
    end
    always @(posedge \clk ) begin
        s96_val_n24 <= s95_val_n24;
    end
    always @(posedge \clk ) begin
        s96_val_n25 <= s95_val_n25;
    end
    always @(posedge \clk ) begin
        s96_val_n26 <= s95_val_n26;
    end
    always @(posedge \clk ) begin
        s96_val_n27 <= s95_val_n27;
    end
    always @(posedge \clk ) begin
        s96_val_n28 <= s95_val_n28;
    end
    always @(posedge \clk ) begin
        s96_val_n29 <= s95_val_n29;
    end
    always @(posedge \clk ) begin
        s96_val_n30 <= s95_val_n30;
    end
    always @(posedge \clk ) begin
        s96_val_n31 <= s95_val_n31;
    end
    always @(posedge \clk ) begin
        s96_val_n32 <= s95_val_n32;
    end
    always @(posedge \clk ) begin
        s96_val_n33 <= s95_val_n33;
    end
    always @(posedge \clk ) begin
        s96_val_n34 <= s95_val_n34;
    end
    always @(posedge \clk ) begin
        s96_val_n35 <= s95_val_n35;
    end
    always @(posedge \clk ) begin
        s96_val_n36 <= s95_val_n36;
    end
    always @(posedge \clk ) begin
        s96_val_n37 <= s95_val_n37;
    end
    always @(posedge \clk ) begin
        s96_val_n38 <= s95_val_n38;
    end
    always @(posedge \clk ) begin
        s96_val_n39 <= s95_val_n39;
    end
    always @(posedge \clk ) begin
        s96_val_n40 <= s95_val_n40;
    end
    always @(posedge \clk ) begin
        s96_val_n41 <= s95_val_n41;
    end
    always @(posedge \clk ) begin
        s96_val_n42 <= s95_val_n42;
    end
    always @(posedge \clk ) begin
        s96_val_n43 <= s95_val_n43;
    end
    always @(posedge \clk ) begin
        s96_val_n44 <= s95_val_n44;
    end
    always @(posedge \clk ) begin
        s96_val_n45 <= s95_val_n45;
    end
    always @(posedge \clk ) begin
        s96_val_n46 <= s95_val_n46;
    end
    always @(posedge \clk ) begin
        \s97_val  <= \s96_val ;
    end
    always @(posedge \clk ) begin
        s97_val_n1 <= s96_val_n1;
    end
    always @(posedge \clk ) begin
        s97_val_n2 <= s96_val_n2;
    end
    always @(posedge \clk ) begin
        s97_val_n3 <= s96_val_n3;
    end
    always @(posedge \clk ) begin
        s97_val_n4 <= s96_val_n4;
    end
    always @(posedge \clk ) begin
        s97_val_n5 <= s96_val_n5;
    end
    always @(posedge \clk ) begin
        s97_val_n6 <= s96_val_n6;
    end
    always @(posedge \clk ) begin
        s97_val_n7 <= s96_val_n7;
    end
    always @(posedge \clk ) begin
        s97_val_n8 <= s96_val_n8;
    end
    always @(posedge \clk ) begin
        s97_val_n9 <= s96_val_n9;
    end
    always @(posedge \clk ) begin
        s97_val_n10 <= s96_val_n10;
    end
    always @(posedge \clk ) begin
        s97_val_n11 <= s96_val_n11;
    end
    always @(posedge \clk ) begin
        s97_val_n12 <= s96_val_n12;
    end
    always @(posedge \clk ) begin
        s97_val_n13 <= s96_val_n13;
    end
    always @(posedge \clk ) begin
        s97_val_n14 <= s96_val_n14;
    end
    always @(posedge \clk ) begin
        s97_val_n15 <= s96_val_n15;
    end
    always @(posedge \clk ) begin
        s97_val_n16 <= s96_val_n16;
    end
    always @(posedge \clk ) begin
        s97_val_n17 <= s96_val_n17;
    end
    always @(posedge \clk ) begin
        s97_val_n18 <= s96_val_n18;
    end
    always @(posedge \clk ) begin
        s97_val_n19 <= s96_val_n19;
    end
    always @(posedge \clk ) begin
        s97_val_n20 <= s96_val_n20;
    end
    always @(posedge \clk ) begin
        s97_val_n21 <= s96_val_n21;
    end
    always @(posedge \clk ) begin
        s97_val_n22 <= s96_val_n22;
    end
    always @(posedge \clk ) begin
        s97_val_n23 <= s96_val_n23;
    end
    always @(posedge \clk ) begin
        s97_val_n24 <= s96_val_n24;
    end
    always @(posedge \clk ) begin
        s97_val_n25 <= s96_val_n25;
    end
    always @(posedge \clk ) begin
        s97_val_n26 <= s96_val_n26;
    end
    always @(posedge \clk ) begin
        s97_val_n27 <= s96_val_n27;
    end
    always @(posedge \clk ) begin
        s97_val_n28 <= s96_val_n28;
    end
    always @(posedge \clk ) begin
        s97_val_n29 <= s96_val_n29;
    end
    always @(posedge \clk ) begin
        s97_val_n30 <= s96_val_n30;
    end
    always @(posedge \clk ) begin
        s97_val_n31 <= s96_val_n31;
    end
    always @(posedge \clk ) begin
        s97_val_n32 <= s96_val_n32;
    end
    always @(posedge \clk ) begin
        s97_val_n33 <= s96_val_n33;
    end
    always @(posedge \clk ) begin
        s97_val_n34 <= s96_val_n34;
    end
    always @(posedge \clk ) begin
        s97_val_n35 <= s96_val_n35;
    end
    always @(posedge \clk ) begin
        s97_val_n36 <= s96_val_n36;
    end
    always @(posedge \clk ) begin
        s97_val_n37 <= s96_val_n37;
    end
    always @(posedge \clk ) begin
        s97_val_n38 <= s96_val_n38;
    end
    always @(posedge \clk ) begin
        s97_val_n39 <= s96_val_n39;
    end
    always @(posedge \clk ) begin
        s97_val_n40 <= s96_val_n40;
    end
    always @(posedge \clk ) begin
        s97_val_n41 <= s96_val_n41;
    end
    always @(posedge \clk ) begin
        s97_val_n42 <= s96_val_n42;
    end
    always @(posedge \clk ) begin
        s97_val_n43 <= s96_val_n43;
    end
    always @(posedge \clk ) begin
        s97_val_n44 <= s96_val_n44;
    end
    always @(posedge \clk ) begin
        s97_val_n45 <= s96_val_n45;
    end
    always @(posedge \clk ) begin
        s97_val_n46 <= s96_val_n46;
    end
    always @(posedge \clk ) begin
        s97_val_n47 <= val_n47;
    end
    always @(posedge \clk ) begin
        \s98_val  <= \s97_val ;
    end
    always @(posedge \clk ) begin
        s98_val_n1 <= s97_val_n1;
    end
    always @(posedge \clk ) begin
        s98_val_n2 <= s97_val_n2;
    end
    always @(posedge \clk ) begin
        s98_val_n3 <= s97_val_n3;
    end
    always @(posedge \clk ) begin
        s98_val_n4 <= s97_val_n4;
    end
    always @(posedge \clk ) begin
        s98_val_n5 <= s97_val_n5;
    end
    always @(posedge \clk ) begin
        s98_val_n6 <= s97_val_n6;
    end
    always @(posedge \clk ) begin
        s98_val_n7 <= s97_val_n7;
    end
    always @(posedge \clk ) begin
        s98_val_n8 <= s97_val_n8;
    end
    always @(posedge \clk ) begin
        s98_val_n9 <= s97_val_n9;
    end
    always @(posedge \clk ) begin
        s98_val_n10 <= s97_val_n10;
    end
    always @(posedge \clk ) begin
        s98_val_n11 <= s97_val_n11;
    end
    always @(posedge \clk ) begin
        s98_val_n12 <= s97_val_n12;
    end
    always @(posedge \clk ) begin
        s98_val_n13 <= s97_val_n13;
    end
    always @(posedge \clk ) begin
        s98_val_n14 <= s97_val_n14;
    end
    always @(posedge \clk ) begin
        s98_val_n15 <= s97_val_n15;
    end
    always @(posedge \clk ) begin
        s98_val_n16 <= s97_val_n16;
    end
    always @(posedge \clk ) begin
        s98_val_n17 <= s97_val_n17;
    end
    always @(posedge \clk ) begin
        s98_val_n18 <= s97_val_n18;
    end
    always @(posedge \clk ) begin
        s98_val_n19 <= s97_val_n19;
    end
    always @(posedge \clk ) begin
        s98_val_n20 <= s97_val_n20;
    end
    always @(posedge \clk ) begin
        s98_val_n21 <= s97_val_n21;
    end
    always @(posedge \clk ) begin
        s98_val_n22 <= s97_val_n22;
    end
    always @(posedge \clk ) begin
        s98_val_n23 <= s97_val_n23;
    end
    always @(posedge \clk ) begin
        s98_val_n24 <= s97_val_n24;
    end
    always @(posedge \clk ) begin
        s98_val_n25 <= s97_val_n25;
    end
    always @(posedge \clk ) begin
        s98_val_n26 <= s97_val_n26;
    end
    always @(posedge \clk ) begin
        s98_val_n27 <= s97_val_n27;
    end
    always @(posedge \clk ) begin
        s98_val_n28 <= s97_val_n28;
    end
    always @(posedge \clk ) begin
        s98_val_n29 <= s97_val_n29;
    end
    always @(posedge \clk ) begin
        s98_val_n30 <= s97_val_n30;
    end
    always @(posedge \clk ) begin
        s98_val_n31 <= s97_val_n31;
    end
    always @(posedge \clk ) begin
        s98_val_n32 <= s97_val_n32;
    end
    always @(posedge \clk ) begin
        s98_val_n33 <= s97_val_n33;
    end
    always @(posedge \clk ) begin
        s98_val_n34 <= s97_val_n34;
    end
    always @(posedge \clk ) begin
        s98_val_n35 <= s97_val_n35;
    end
    always @(posedge \clk ) begin
        s98_val_n36 <= s97_val_n36;
    end
    always @(posedge \clk ) begin
        s98_val_n37 <= s97_val_n37;
    end
    always @(posedge \clk ) begin
        s98_val_n38 <= s97_val_n38;
    end
    always @(posedge \clk ) begin
        s98_val_n39 <= s97_val_n39;
    end
    always @(posedge \clk ) begin
        s98_val_n40 <= s97_val_n40;
    end
    always @(posedge \clk ) begin
        s98_val_n41 <= s97_val_n41;
    end
    always @(posedge \clk ) begin
        s98_val_n42 <= s97_val_n42;
    end
    always @(posedge \clk ) begin
        s98_val_n43 <= s97_val_n43;
    end
    always @(posedge \clk ) begin
        s98_val_n44 <= s97_val_n44;
    end
    always @(posedge \clk ) begin
        s98_val_n45 <= s97_val_n45;
    end
    always @(posedge \clk ) begin
        s98_val_n46 <= s97_val_n46;
    end
    always @(posedge \clk ) begin
        s98_val_n47 <= s97_val_n47;
    end
    always @(posedge \clk ) begin
        \s99_val  <= \s98_val ;
    end
    always @(posedge \clk ) begin
        s99_val_n1 <= s98_val_n1;
    end
    always @(posedge \clk ) begin
        s99_val_n2 <= s98_val_n2;
    end
    always @(posedge \clk ) begin
        s99_val_n3 <= s98_val_n3;
    end
    always @(posedge \clk ) begin
        s99_val_n4 <= s98_val_n4;
    end
    always @(posedge \clk ) begin
        s99_val_n5 <= s98_val_n5;
    end
    always @(posedge \clk ) begin
        s99_val_n6 <= s98_val_n6;
    end
    always @(posedge \clk ) begin
        s99_val_n7 <= s98_val_n7;
    end
    always @(posedge \clk ) begin
        s99_val_n8 <= s98_val_n8;
    end
    always @(posedge \clk ) begin
        s99_val_n9 <= s98_val_n9;
    end
    always @(posedge \clk ) begin
        s99_val_n10 <= s98_val_n10;
    end
    always @(posedge \clk ) begin
        s99_val_n11 <= s98_val_n11;
    end
    always @(posedge \clk ) begin
        s99_val_n12 <= s98_val_n12;
    end
    always @(posedge \clk ) begin
        s99_val_n13 <= s98_val_n13;
    end
    always @(posedge \clk ) begin
        s99_val_n14 <= s98_val_n14;
    end
    always @(posedge \clk ) begin
        s99_val_n15 <= s98_val_n15;
    end
    always @(posedge \clk ) begin
        s99_val_n16 <= s98_val_n16;
    end
    always @(posedge \clk ) begin
        s99_val_n17 <= s98_val_n17;
    end
    always @(posedge \clk ) begin
        s99_val_n18 <= s98_val_n18;
    end
    always @(posedge \clk ) begin
        s99_val_n19 <= s98_val_n19;
    end
    always @(posedge \clk ) begin
        s99_val_n20 <= s98_val_n20;
    end
    always @(posedge \clk ) begin
        s99_val_n21 <= s98_val_n21;
    end
    always @(posedge \clk ) begin
        s99_val_n22 <= s98_val_n22;
    end
    always @(posedge \clk ) begin
        s99_val_n23 <= s98_val_n23;
    end
    always @(posedge \clk ) begin
        s99_val_n24 <= s98_val_n24;
    end
    always @(posedge \clk ) begin
        s99_val_n25 <= s98_val_n25;
    end
    always @(posedge \clk ) begin
        s99_val_n26 <= s98_val_n26;
    end
    always @(posedge \clk ) begin
        s99_val_n27 <= s98_val_n27;
    end
    always @(posedge \clk ) begin
        s99_val_n28 <= s98_val_n28;
    end
    always @(posedge \clk ) begin
        s99_val_n29 <= s98_val_n29;
    end
    always @(posedge \clk ) begin
        s99_val_n30 <= s98_val_n30;
    end
    always @(posedge \clk ) begin
        s99_val_n31 <= s98_val_n31;
    end
    always @(posedge \clk ) begin
        s99_val_n32 <= s98_val_n32;
    end
    always @(posedge \clk ) begin
        s99_val_n33 <= s98_val_n33;
    end
    always @(posedge \clk ) begin
        s99_val_n34 <= s98_val_n34;
    end
    always @(posedge \clk ) begin
        s99_val_n35 <= s98_val_n35;
    end
    always @(posedge \clk ) begin
        s99_val_n36 <= s98_val_n36;
    end
    always @(posedge \clk ) begin
        s99_val_n37 <= s98_val_n37;
    end
    always @(posedge \clk ) begin
        s99_val_n38 <= s98_val_n38;
    end
    always @(posedge \clk ) begin
        s99_val_n39 <= s98_val_n39;
    end
    always @(posedge \clk ) begin
        s99_val_n40 <= s98_val_n40;
    end
    always @(posedge \clk ) begin
        s99_val_n41 <= s98_val_n41;
    end
    always @(posedge \clk ) begin
        s99_val_n42 <= s98_val_n42;
    end
    always @(posedge \clk ) begin
        s99_val_n43 <= s98_val_n43;
    end
    always @(posedge \clk ) begin
        s99_val_n44 <= s98_val_n44;
    end
    always @(posedge \clk ) begin
        s99_val_n45 <= s98_val_n45;
    end
    always @(posedge \clk ) begin
        s99_val_n46 <= s98_val_n46;
    end
    always @(posedge \clk ) begin
        s99_val_n47 <= s98_val_n47;
    end
    always @(posedge \clk ) begin
        s99_val_n48 <= val_n48;
    end
    always @(posedge \clk ) begin
        \s100_val  <= \s99_val ;
    end
    always @(posedge \clk ) begin
        s100_val_n1 <= s99_val_n1;
    end
    always @(posedge \clk ) begin
        s100_val_n2 <= s99_val_n2;
    end
    always @(posedge \clk ) begin
        s100_val_n3 <= s99_val_n3;
    end
    always @(posedge \clk ) begin
        s100_val_n4 <= s99_val_n4;
    end
    always @(posedge \clk ) begin
        s100_val_n5 <= s99_val_n5;
    end
    always @(posedge \clk ) begin
        s100_val_n6 <= s99_val_n6;
    end
    always @(posedge \clk ) begin
        s100_val_n7 <= s99_val_n7;
    end
    always @(posedge \clk ) begin
        s100_val_n8 <= s99_val_n8;
    end
    always @(posedge \clk ) begin
        s100_val_n9 <= s99_val_n9;
    end
    always @(posedge \clk ) begin
        s100_val_n10 <= s99_val_n10;
    end
    always @(posedge \clk ) begin
        s100_val_n11 <= s99_val_n11;
    end
    always @(posedge \clk ) begin
        s100_val_n12 <= s99_val_n12;
    end
    always @(posedge \clk ) begin
        s100_val_n13 <= s99_val_n13;
    end
    always @(posedge \clk ) begin
        s100_val_n14 <= s99_val_n14;
    end
    always @(posedge \clk ) begin
        s100_val_n15 <= s99_val_n15;
    end
    always @(posedge \clk ) begin
        s100_val_n16 <= s99_val_n16;
    end
    always @(posedge \clk ) begin
        s100_val_n17 <= s99_val_n17;
    end
    always @(posedge \clk ) begin
        s100_val_n18 <= s99_val_n18;
    end
    always @(posedge \clk ) begin
        s100_val_n19 <= s99_val_n19;
    end
    always @(posedge \clk ) begin
        s100_val_n20 <= s99_val_n20;
    end
    always @(posedge \clk ) begin
        s100_val_n21 <= s99_val_n21;
    end
    always @(posedge \clk ) begin
        s100_val_n22 <= s99_val_n22;
    end
    always @(posedge \clk ) begin
        s100_val_n23 <= s99_val_n23;
    end
    always @(posedge \clk ) begin
        s100_val_n24 <= s99_val_n24;
    end
    always @(posedge \clk ) begin
        s100_val_n25 <= s99_val_n25;
    end
    always @(posedge \clk ) begin
        s100_val_n26 <= s99_val_n26;
    end
    always @(posedge \clk ) begin
        s100_val_n27 <= s99_val_n27;
    end
    always @(posedge \clk ) begin
        s100_val_n28 <= s99_val_n28;
    end
    always @(posedge \clk ) begin
        s100_val_n29 <= s99_val_n29;
    end
    always @(posedge \clk ) begin
        s100_val_n30 <= s99_val_n30;
    end
    always @(posedge \clk ) begin
        s100_val_n31 <= s99_val_n31;
    end
    always @(posedge \clk ) begin
        s100_val_n32 <= s99_val_n32;
    end
    always @(posedge \clk ) begin
        s100_val_n33 <= s99_val_n33;
    end
    always @(posedge \clk ) begin
        s100_val_n34 <= s99_val_n34;
    end
    always @(posedge \clk ) begin
        s100_val_n35 <= s99_val_n35;
    end
    always @(posedge \clk ) begin
        s100_val_n36 <= s99_val_n36;
    end
    always @(posedge \clk ) begin
        s100_val_n37 <= s99_val_n37;
    end
    always @(posedge \clk ) begin
        s100_val_n38 <= s99_val_n38;
    end
    always @(posedge \clk ) begin
        s100_val_n39 <= s99_val_n39;
    end
    always @(posedge \clk ) begin
        s100_val_n40 <= s99_val_n40;
    end
    always @(posedge \clk ) begin
        s100_val_n41 <= s99_val_n41;
    end
    always @(posedge \clk ) begin
        s100_val_n42 <= s99_val_n42;
    end
    always @(posedge \clk ) begin
        s100_val_n43 <= s99_val_n43;
    end
    always @(posedge \clk ) begin
        s100_val_n44 <= s99_val_n44;
    end
    always @(posedge \clk ) begin
        s100_val_n45 <= s99_val_n45;
    end
    always @(posedge \clk ) begin
        s100_val_n46 <= s99_val_n46;
    end
    always @(posedge \clk ) begin
        s100_val_n47 <= s99_val_n47;
    end
    always @(posedge \clk ) begin
        s100_val_n48 <= s99_val_n48;
    end
    (* src = "src/sreg.spade:25,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_0(.clk_i(\clk ), .val_i(\s2_val ), .output__(val_n1));
    (* src = "src/sreg.spade:27,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_1(.clk_i(\clk ), .val_i(val_n1), .output__(val_n2));
    (* src = "src/sreg.spade:29,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_2(.clk_i(\clk ), .val_i(val_n2), .output__(val_n3));
    (* src = "src/sreg.spade:31,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_3(.clk_i(\clk ), .val_i(val_n3), .output__(val_n4));
    (* src = "src/sreg.spade:33,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_4(.clk_i(\clk ), .val_i(val_n4), .output__(val_n5));
    (* src = "src/sreg.spade:35,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_5(.clk_i(\clk ), .val_i(val_n5), .output__(val_n6));
    (* src = "src/sreg.spade:37,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_6(.clk_i(\clk ), .val_i(val_n6), .output__(val_n7));
    (* src = "src/sreg.spade:39,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_7(.clk_i(\clk ), .val_i(val_n7), .output__(val_n8));
    (* src = "src/sreg.spade:41,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_8(.clk_i(\clk ), .val_i(val_n8), .output__(val_n9));
    (* src = "src/sreg.spade:43,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_9(.clk_i(\clk ), .val_i(val_n9), .output__(val_n10));
    (* src = "src/sreg.spade:45,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_10(.clk_i(\clk ), .val_i(val_n10), .output__(val_n11));
    (* src = "src/sreg.spade:47,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_11(.clk_i(\clk ), .val_i(val_n11), .output__(val_n12));
    (* src = "src/sreg.spade:49,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_12(.clk_i(\clk ), .val_i(val_n12), .output__(val_n13));
    (* src = "src/sreg.spade:51,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_13(.clk_i(\clk ), .val_i(val_n13), .output__(val_n14));
    (* src = "src/sreg.spade:53,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_14(.clk_i(\clk ), .val_i(val_n14), .output__(val_n15));
    (* src = "src/sreg.spade:55,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_15(.clk_i(\clk ), .val_i(val_n15), .output__(val_n16));
    (* src = "src/sreg.spade:57,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_16(.clk_i(\clk ), .val_i(val_n16), .output__(val_n17));
    (* src = "src/sreg.spade:59,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_17(.clk_i(\clk ), .val_i(val_n17), .output__(val_n18));
    (* src = "src/sreg.spade:61,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_18(.clk_i(\clk ), .val_i(val_n18), .output__(val_n19));
    (* src = "src/sreg.spade:63,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_19(.clk_i(\clk ), .val_i(val_n19), .output__(val_n20));
    (* src = "src/sreg.spade:65,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_20(.clk_i(\clk ), .val_i(val_n20), .output__(val_n21));
    (* src = "src/sreg.spade:67,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_21(.clk_i(\clk ), .val_i(val_n21), .output__(val_n22));
    (* src = "src/sreg.spade:69,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_22(.clk_i(\clk ), .val_i(val_n22), .output__(val_n23));
    (* src = "src/sreg.spade:71,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_23(.clk_i(\clk ), .val_i(val_n23), .output__(val_n24));
    (* src = "src/sreg.spade:73,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_24(.clk_i(\clk ), .val_i(val_n24), .output__(val_n25));
    (* src = "src/sreg.spade:75,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_25(.clk_i(\clk ), .val_i(val_n25), .output__(val_n26));
    (* src = "src/sreg.spade:77,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_26(.clk_i(\clk ), .val_i(val_n26), .output__(val_n27));
    (* src = "src/sreg.spade:79,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_27(.clk_i(\clk ), .val_i(val_n27), .output__(val_n28));
    (* src = "src/sreg.spade:81,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_28(.clk_i(\clk ), .val_i(val_n28), .output__(val_n29));
    (* src = "src/sreg.spade:83,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_29(.clk_i(\clk ), .val_i(val_n29), .output__(val_n30));
    (* src = "src/sreg.spade:85,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_30(.clk_i(\clk ), .val_i(val_n30), .output__(val_n31));
    (* src = "src/sreg.spade:87,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_31(.clk_i(\clk ), .val_i(val_n31), .output__(val_n32));
    (* src = "src/sreg.spade:89,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_32(.clk_i(\clk ), .val_i(val_n32), .output__(val_n33));
    (* src = "src/sreg.spade:91,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_33(.clk_i(\clk ), .val_i(val_n33), .output__(val_n34));
    (* src = "src/sreg.spade:93,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_34(.clk_i(\clk ), .val_i(val_n34), .output__(val_n35));
    (* src = "src/sreg.spade:95,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_35(.clk_i(\clk ), .val_i(val_n35), .output__(val_n36));
    (* src = "src/sreg.spade:97,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_36(.clk_i(\clk ), .val_i(val_n36), .output__(val_n37));
    (* src = "src/sreg.spade:99,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_37(.clk_i(\clk ), .val_i(val_n37), .output__(val_n38));
    (* src = "src/sreg.spade:101,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_38(.clk_i(\clk ), .val_i(val_n38), .output__(val_n39));
    (* src = "src/sreg.spade:103,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_39(.clk_i(\clk ), .val_i(val_n39), .output__(val_n40));
    (* src = "src/sreg.spade:105,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_40(.clk_i(\clk ), .val_i(val_n40), .output__(val_n41));
    (* src = "src/sreg.spade:107,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_41(.clk_i(\clk ), .val_i(val_n41), .output__(val_n42));
    (* src = "src/sreg.spade:109,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_42(.clk_i(\clk ), .val_i(val_n42), .output__(val_n43));
    (* src = "src/sreg.spade:111,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_43(.clk_i(\clk ), .val_i(val_n43), .output__(val_n44));
    (* src = "src/sreg.spade:113,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_44(.clk_i(\clk ), .val_i(val_n44), .output__(val_n45));
    (* src = "src/sreg.spade:115,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_45(.clk_i(\clk ), .val_i(val_n45), .output__(val_n46));
    (* src = "src/sreg.spade:117,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_46(.clk_i(\clk ), .val_i(val_n46), .output__(val_n47));
    (* src = "src/sreg.spade:119,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_47(.clk_i(\clk ), .val_i(val_n47), .output__(val_n48));
    (* src = "src/sreg.spade:121,19" *)
    \tt07_delay_line_tmng::sreg::inv_reg  inv_reg_48(.clk_i(\clk ), .val_i(val_n48), .output__(val_n49));
    assign output__ = val_n49;
endmodule

module \tt07_delay_line_tmng::sreg::shift_reg  (
        input clk_i,
        input val_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "tt07_delay_line_tmng::sreg::shift_reg" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \tt07_delay_line_tmng::sreg::shift_reg );
        end
    end
    `endif
    logic \clk ;
    assign \clk  = clk_i;
    logic \val ;
    assign \val  = val_i;
    (* src = "src/sreg.spade:128,5" *)
    reg \s1_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s2_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s3_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s4_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s5_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s6_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s7_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s8_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s9_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s10_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s11_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s12_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s13_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s14_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s15_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s16_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s17_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s18_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s19_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s20_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s21_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s22_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s23_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s24_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s25_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s26_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s27_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s28_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s29_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s30_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s31_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s32_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s33_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s34_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s35_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s36_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s37_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s38_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s39_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s40_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s41_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s42_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s43_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s44_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s45_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s46_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s47_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s48_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s49_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s50_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s51_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s52_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s53_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s54_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s55_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s56_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s57_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s58_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s59_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s60_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s61_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s62_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s63_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s64_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s65_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s66_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s67_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s68_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s69_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s70_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s71_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s72_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s73_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s74_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s75_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s76_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s77_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s78_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s79_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s80_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s81_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s82_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s83_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s84_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s85_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s86_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s87_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s88_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s89_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s90_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s91_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s92_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s93_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s94_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s95_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s96_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s97_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s98_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s99_val ;
    (* src = "src/sreg.spade:128,5" *)
    reg \s100_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg \s101_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s101_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s102_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s102_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s103_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s103_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s104_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s104_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s105_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s105_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s106_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s106_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s107_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s107_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s108_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s108_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s109_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s109_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s110_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s110_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s111_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s111_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s112_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s112_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s113_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s113_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s114_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s114_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s115_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s115_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s116_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s116_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s117_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s117_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s118_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s118_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s119_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s119_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s120_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s120_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s121_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s121_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s122_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s122_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s123_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s123_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s124_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s124_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s125_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s125_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s126_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s126_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s127_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s127_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s128_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s128_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s129_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s129_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s130_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s130_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s131_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s131_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s132_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s132_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s133_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s133_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s134_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s134_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s135_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s135_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s136_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s136_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s137_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s137_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s138_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s138_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s139_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s139_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s140_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s140_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s141_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s141_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s142_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s142_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s143_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s143_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s144_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s144_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s145_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s145_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s146_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s146_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s147_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s147_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s148_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s148_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s149_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s149_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s150_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s150_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s151_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s151_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s152_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s152_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s153_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s153_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s154_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s154_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s155_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s155_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s156_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s156_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s157_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s157_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s158_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s158_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s159_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s159_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s160_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s160_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s161_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s161_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s162_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s162_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s163_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s163_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s164_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s164_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s165_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s165_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s166_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s166_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s167_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s167_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s168_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s168_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s169_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s169_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s170_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s170_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s171_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s171_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s172_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s172_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s173_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s173_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s174_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s174_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s175_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s175_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s176_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s176_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s177_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s177_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s178_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s178_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s179_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s179_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s180_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s180_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s181_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s181_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s182_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s182_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s183_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s183_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s184_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s184_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s185_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s185_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s186_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s186_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s187_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s187_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s188_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s188_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s189_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s189_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s190_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s190_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s191_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s191_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s192_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s192_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s193_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s193_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s194_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s194_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s195_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s195_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s196_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s196_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s197_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s197_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s198_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s198_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s199_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s199_val_n1;
    (* src = "src/sreg.spade:130,5" *)
    reg \s200_val ;
    (* src = "src/sreg.spade:130,5" *)
    reg s200_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg \s201_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s201_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s201_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s202_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s202_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s202_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s203_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s203_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s203_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s204_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s204_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s204_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s205_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s205_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s205_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s206_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s206_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s206_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s207_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s207_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s207_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s208_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s208_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s208_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s209_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s209_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s209_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s210_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s210_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s210_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s211_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s211_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s211_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s212_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s212_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s212_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s213_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s213_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s213_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s214_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s214_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s214_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s215_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s215_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s215_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s216_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s216_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s216_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s217_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s217_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s217_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s218_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s218_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s218_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s219_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s219_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s219_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s220_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s220_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s220_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s221_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s221_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s221_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s222_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s222_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s222_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s223_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s223_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s223_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s224_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s224_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s224_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s225_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s225_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s225_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s226_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s226_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s226_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s227_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s227_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s227_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s228_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s228_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s228_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s229_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s229_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s229_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s230_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s230_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s230_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s231_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s231_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s231_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s232_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s232_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s232_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s233_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s233_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s233_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s234_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s234_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s234_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s235_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s235_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s235_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s236_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s236_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s236_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s237_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s237_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s237_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s238_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s238_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s238_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s239_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s239_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s239_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s240_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s240_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s240_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s241_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s241_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s241_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s242_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s242_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s242_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s243_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s243_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s243_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s244_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s244_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s244_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s245_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s245_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s245_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s246_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s246_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s246_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s247_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s247_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s247_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s248_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s248_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s248_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s249_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s249_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s249_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s250_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s250_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s250_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s251_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s251_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s251_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s252_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s252_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s252_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s253_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s253_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s253_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s254_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s254_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s254_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s255_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s255_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s255_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s256_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s256_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s256_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s257_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s257_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s257_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s258_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s258_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s258_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s259_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s259_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s259_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s260_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s260_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s260_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s261_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s261_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s261_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s262_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s262_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s262_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s263_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s263_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s263_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s264_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s264_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s264_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s265_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s265_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s265_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s266_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s266_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s266_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s267_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s267_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s267_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s268_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s268_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s268_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s269_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s269_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s269_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s270_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s270_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s270_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s271_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s271_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s271_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s272_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s272_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s272_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s273_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s273_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s273_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s274_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s274_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s274_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s275_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s275_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s275_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s276_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s276_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s276_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s277_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s277_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s277_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s278_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s278_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s278_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s279_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s279_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s279_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s280_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s280_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s280_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s281_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s281_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s281_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s282_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s282_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s282_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s283_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s283_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s283_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s284_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s284_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s284_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s285_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s285_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s285_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s286_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s286_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s286_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s287_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s287_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s287_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s288_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s288_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s288_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s289_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s289_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s289_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s290_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s290_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s290_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s291_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s291_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s291_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s292_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s292_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s292_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s293_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s293_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s293_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s294_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s294_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s294_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s295_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s295_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s295_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s296_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s296_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s296_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s297_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s297_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s297_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s298_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s298_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s298_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s299_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s299_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s299_val_n2;
    (* src = "src/sreg.spade:132,5" *)
    reg \s300_val ;
    (* src = "src/sreg.spade:132,5" *)
    reg s300_val_n1;
    (* src = "src/sreg.spade:132,5" *)
    reg s300_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg \s301_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s301_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s301_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s301_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s302_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s302_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s302_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s302_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s303_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s303_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s303_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s303_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s304_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s304_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s304_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s304_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s305_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s305_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s305_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s305_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s306_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s306_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s306_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s306_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s307_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s307_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s307_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s307_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s308_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s308_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s308_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s308_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s309_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s309_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s309_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s309_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s310_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s310_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s310_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s310_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s311_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s311_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s311_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s311_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s312_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s312_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s312_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s312_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s313_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s313_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s313_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s313_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s314_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s314_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s314_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s314_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s315_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s315_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s315_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s315_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s316_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s316_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s316_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s316_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s317_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s317_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s317_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s317_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s318_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s318_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s318_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s318_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s319_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s319_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s319_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s319_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s320_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s320_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s320_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s320_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s321_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s321_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s321_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s321_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s322_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s322_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s322_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s322_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s323_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s323_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s323_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s323_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s324_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s324_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s324_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s324_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s325_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s325_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s325_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s325_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s326_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s326_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s326_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s326_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s327_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s327_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s327_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s327_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s328_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s328_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s328_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s328_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s329_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s329_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s329_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s329_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s330_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s330_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s330_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s330_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s331_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s331_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s331_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s331_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s332_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s332_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s332_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s332_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s333_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s333_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s333_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s333_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s334_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s334_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s334_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s334_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s335_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s335_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s335_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s335_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s336_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s336_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s336_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s336_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s337_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s337_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s337_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s337_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s338_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s338_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s338_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s338_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s339_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s339_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s339_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s339_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s340_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s340_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s340_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s340_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s341_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s341_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s341_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s341_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s342_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s342_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s342_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s342_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s343_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s343_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s343_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s343_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s344_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s344_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s344_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s344_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s345_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s345_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s345_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s345_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s346_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s346_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s346_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s346_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s347_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s347_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s347_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s347_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s348_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s348_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s348_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s348_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s349_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s349_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s349_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s349_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s350_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s350_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s350_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s350_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s351_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s351_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s351_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s351_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s352_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s352_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s352_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s352_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s353_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s353_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s353_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s353_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s354_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s354_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s354_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s354_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s355_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s355_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s355_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s355_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s356_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s356_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s356_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s356_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s357_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s357_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s357_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s357_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s358_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s358_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s358_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s358_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s359_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s359_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s359_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s359_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s360_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s360_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s360_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s360_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s361_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s361_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s361_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s361_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s362_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s362_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s362_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s362_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s363_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s363_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s363_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s363_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s364_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s364_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s364_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s364_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s365_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s365_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s365_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s365_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s366_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s366_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s366_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s366_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s367_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s367_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s367_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s367_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s368_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s368_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s368_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s368_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s369_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s369_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s369_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s369_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s370_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s370_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s370_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s370_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s371_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s371_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s371_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s371_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s372_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s372_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s372_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s372_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s373_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s373_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s373_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s373_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s374_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s374_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s374_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s374_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s375_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s375_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s375_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s375_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s376_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s376_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s376_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s376_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s377_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s377_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s377_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s377_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s378_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s378_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s378_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s378_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s379_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s379_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s379_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s379_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s380_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s380_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s380_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s380_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s381_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s381_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s381_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s381_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s382_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s382_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s382_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s382_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s383_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s383_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s383_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s383_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s384_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s384_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s384_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s384_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s385_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s385_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s385_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s385_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s386_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s386_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s386_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s386_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s387_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s387_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s387_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s387_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s388_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s388_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s388_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s388_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s389_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s389_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s389_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s389_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s390_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s390_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s390_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s390_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s391_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s391_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s391_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s391_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s392_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s392_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s392_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s392_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s393_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s393_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s393_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s393_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s394_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s394_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s394_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s394_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s395_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s395_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s395_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s395_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s396_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s396_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s396_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s396_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s397_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s397_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s397_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s397_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s398_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s398_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s398_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s398_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s399_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s399_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s399_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s399_val_n3;
    (* src = "src/sreg.spade:134,5" *)
    reg \s400_val ;
    (* src = "src/sreg.spade:134,5" *)
    reg s400_val_n1;
    (* src = "src/sreg.spade:134,5" *)
    reg s400_val_n2;
    (* src = "src/sreg.spade:134,5" *)
    reg s400_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg \s401_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s401_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s401_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s401_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s401_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s402_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s402_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s402_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s402_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s402_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s403_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s403_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s403_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s403_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s403_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s404_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s404_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s404_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s404_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s404_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s405_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s405_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s405_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s405_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s405_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s406_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s406_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s406_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s406_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s406_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s407_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s407_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s407_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s407_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s407_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s408_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s408_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s408_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s408_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s408_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s409_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s409_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s409_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s409_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s409_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s410_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s410_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s410_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s410_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s410_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s411_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s411_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s411_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s411_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s411_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s412_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s412_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s412_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s412_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s412_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s413_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s413_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s413_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s413_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s413_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s414_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s414_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s414_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s414_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s414_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s415_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s415_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s415_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s415_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s415_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s416_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s416_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s416_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s416_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s416_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s417_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s417_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s417_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s417_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s417_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s418_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s418_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s418_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s418_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s418_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s419_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s419_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s419_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s419_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s419_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s420_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s420_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s420_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s420_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s420_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s421_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s421_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s421_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s421_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s421_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s422_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s422_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s422_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s422_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s422_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s423_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s423_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s423_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s423_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s423_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s424_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s424_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s424_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s424_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s424_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s425_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s425_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s425_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s425_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s425_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s426_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s426_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s426_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s426_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s426_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s427_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s427_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s427_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s427_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s427_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s428_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s428_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s428_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s428_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s428_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s429_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s429_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s429_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s429_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s429_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s430_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s430_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s430_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s430_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s430_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s431_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s431_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s431_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s431_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s431_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s432_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s432_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s432_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s432_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s432_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s433_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s433_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s433_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s433_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s433_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s434_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s434_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s434_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s434_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s434_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s435_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s435_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s435_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s435_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s435_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s436_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s436_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s436_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s436_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s436_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s437_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s437_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s437_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s437_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s437_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s438_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s438_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s438_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s438_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s438_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s439_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s439_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s439_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s439_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s439_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s440_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s440_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s440_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s440_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s440_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s441_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s441_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s441_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s441_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s441_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s442_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s442_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s442_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s442_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s442_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s443_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s443_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s443_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s443_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s443_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s444_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s444_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s444_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s444_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s444_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s445_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s445_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s445_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s445_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s445_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s446_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s446_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s446_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s446_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s446_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s447_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s447_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s447_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s447_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s447_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s448_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s448_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s448_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s448_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s448_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s449_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s449_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s449_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s449_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s449_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s450_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s450_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s450_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s450_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s450_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s451_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s451_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s451_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s451_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s451_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s452_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s452_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s452_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s452_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s452_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s453_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s453_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s453_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s453_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s453_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s454_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s454_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s454_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s454_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s454_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s455_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s455_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s455_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s455_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s455_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s456_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s456_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s456_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s456_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s456_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s457_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s457_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s457_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s457_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s457_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s458_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s458_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s458_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s458_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s458_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s459_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s459_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s459_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s459_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s459_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s460_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s460_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s460_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s460_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s460_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s461_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s461_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s461_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s461_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s461_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s462_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s462_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s462_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s462_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s462_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s463_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s463_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s463_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s463_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s463_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s464_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s464_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s464_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s464_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s464_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s465_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s465_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s465_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s465_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s465_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s466_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s466_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s466_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s466_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s466_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s467_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s467_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s467_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s467_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s467_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s468_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s468_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s468_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s468_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s468_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s469_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s469_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s469_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s469_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s469_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s470_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s470_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s470_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s470_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s470_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s471_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s471_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s471_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s471_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s471_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s472_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s472_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s472_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s472_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s472_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s473_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s473_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s473_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s473_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s473_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s474_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s474_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s474_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s474_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s474_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s475_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s475_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s475_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s475_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s475_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s476_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s476_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s476_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s476_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s476_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s477_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s477_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s477_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s477_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s477_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s478_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s478_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s478_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s478_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s478_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s479_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s479_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s479_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s479_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s479_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s480_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s480_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s480_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s480_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s480_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s481_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s481_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s481_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s481_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s481_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s482_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s482_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s482_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s482_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s482_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s483_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s483_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s483_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s483_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s483_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s484_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s484_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s484_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s484_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s484_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s485_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s485_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s485_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s485_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s485_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s486_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s486_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s486_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s486_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s486_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s487_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s487_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s487_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s487_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s487_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s488_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s488_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s488_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s488_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s488_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s489_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s489_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s489_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s489_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s489_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s490_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s490_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s490_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s490_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s490_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s491_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s491_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s491_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s491_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s491_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s492_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s492_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s492_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s492_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s492_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s493_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s493_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s493_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s493_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s493_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s494_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s494_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s494_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s494_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s494_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s495_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s495_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s495_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s495_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s495_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s496_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s496_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s496_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s496_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s496_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s497_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s497_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s497_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s497_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s497_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s498_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s498_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s498_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s498_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s498_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s499_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s499_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s499_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s499_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s499_val_n4;
    (* src = "src/sreg.spade:136,5" *)
    reg \s500_val ;
    (* src = "src/sreg.spade:136,5" *)
    reg s500_val_n1;
    (* src = "src/sreg.spade:136,5" *)
    reg s500_val_n2;
    (* src = "src/sreg.spade:136,5" *)
    reg s500_val_n3;
    (* src = "src/sreg.spade:136,5" *)
    reg s500_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg \s501_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s501_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s501_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s501_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s501_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s501_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s502_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s502_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s502_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s502_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s502_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s502_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s503_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s503_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s503_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s503_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s503_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s503_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s504_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s504_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s504_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s504_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s504_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s504_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s505_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s505_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s505_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s505_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s505_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s505_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s506_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s506_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s506_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s506_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s506_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s506_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s507_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s507_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s507_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s507_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s507_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s507_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s508_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s508_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s508_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s508_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s508_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s508_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s509_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s509_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s509_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s509_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s509_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s509_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s510_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s510_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s510_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s510_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s510_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s510_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s511_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s511_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s511_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s511_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s511_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s511_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s512_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s512_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s512_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s512_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s512_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s512_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s513_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s513_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s513_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s513_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s513_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s513_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s514_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s514_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s514_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s514_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s514_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s514_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s515_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s515_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s515_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s515_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s515_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s515_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s516_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s516_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s516_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s516_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s516_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s516_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s517_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s517_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s517_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s517_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s517_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s517_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s518_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s518_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s518_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s518_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s518_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s518_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s519_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s519_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s519_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s519_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s519_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s519_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s520_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s520_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s520_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s520_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s520_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s520_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s521_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s521_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s521_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s521_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s521_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s521_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s522_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s522_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s522_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s522_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s522_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s522_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s523_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s523_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s523_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s523_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s523_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s523_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s524_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s524_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s524_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s524_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s524_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s524_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s525_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s525_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s525_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s525_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s525_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s525_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s526_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s526_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s526_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s526_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s526_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s526_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s527_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s527_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s527_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s527_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s527_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s527_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s528_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s528_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s528_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s528_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s528_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s528_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s529_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s529_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s529_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s529_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s529_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s529_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s530_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s530_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s530_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s530_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s530_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s530_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s531_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s531_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s531_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s531_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s531_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s531_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s532_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s532_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s532_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s532_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s532_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s532_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s533_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s533_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s533_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s533_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s533_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s533_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s534_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s534_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s534_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s534_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s534_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s534_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s535_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s535_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s535_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s535_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s535_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s535_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s536_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s536_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s536_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s536_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s536_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s536_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s537_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s537_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s537_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s537_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s537_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s537_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s538_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s538_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s538_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s538_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s538_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s538_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s539_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s539_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s539_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s539_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s539_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s539_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s540_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s540_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s540_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s540_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s540_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s540_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s541_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s541_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s541_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s541_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s541_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s541_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s542_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s542_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s542_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s542_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s542_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s542_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s543_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s543_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s543_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s543_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s543_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s543_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s544_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s544_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s544_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s544_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s544_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s544_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s545_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s545_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s545_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s545_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s545_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s545_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s546_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s546_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s546_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s546_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s546_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s546_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s547_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s547_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s547_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s547_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s547_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s547_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s548_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s548_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s548_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s548_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s548_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s548_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s549_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s549_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s549_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s549_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s549_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s549_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s550_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s550_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s550_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s550_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s550_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s550_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s551_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s551_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s551_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s551_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s551_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s551_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s552_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s552_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s552_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s552_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s552_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s552_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s553_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s553_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s553_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s553_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s553_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s553_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s554_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s554_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s554_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s554_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s554_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s554_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s555_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s555_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s555_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s555_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s555_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s555_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s556_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s556_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s556_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s556_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s556_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s556_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s557_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s557_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s557_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s557_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s557_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s557_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s558_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s558_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s558_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s558_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s558_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s558_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s559_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s559_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s559_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s559_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s559_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s559_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s560_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s560_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s560_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s560_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s560_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s560_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s561_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s561_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s561_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s561_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s561_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s561_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s562_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s562_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s562_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s562_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s562_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s562_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s563_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s563_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s563_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s563_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s563_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s563_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s564_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s564_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s564_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s564_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s564_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s564_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s565_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s565_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s565_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s565_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s565_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s565_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s566_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s566_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s566_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s566_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s566_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s566_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s567_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s567_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s567_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s567_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s567_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s567_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s568_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s568_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s568_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s568_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s568_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s568_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s569_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s569_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s569_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s569_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s569_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s569_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s570_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s570_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s570_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s570_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s570_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s570_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s571_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s571_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s571_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s571_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s571_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s571_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s572_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s572_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s572_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s572_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s572_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s572_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s573_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s573_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s573_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s573_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s573_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s573_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s574_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s574_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s574_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s574_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s574_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s574_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s575_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s575_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s575_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s575_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s575_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s575_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s576_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s576_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s576_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s576_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s576_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s576_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s577_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s577_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s577_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s577_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s577_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s577_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s578_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s578_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s578_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s578_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s578_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s578_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s579_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s579_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s579_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s579_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s579_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s579_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s580_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s580_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s580_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s580_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s580_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s580_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s581_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s581_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s581_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s581_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s581_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s581_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s582_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s582_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s582_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s582_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s582_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s582_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s583_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s583_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s583_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s583_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s583_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s583_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s584_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s584_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s584_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s584_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s584_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s584_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s585_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s585_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s585_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s585_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s585_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s585_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s586_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s586_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s586_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s586_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s586_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s586_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s587_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s587_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s587_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s587_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s587_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s587_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s588_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s588_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s588_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s588_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s588_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s588_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s589_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s589_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s589_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s589_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s589_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s589_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s590_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s590_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s590_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s590_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s590_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s590_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s591_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s591_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s591_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s591_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s591_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s591_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s592_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s592_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s592_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s592_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s592_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s592_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s593_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s593_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s593_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s593_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s593_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s593_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s594_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s594_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s594_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s594_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s594_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s594_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s595_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s595_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s595_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s595_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s595_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s595_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s596_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s596_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s596_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s596_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s596_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s596_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s597_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s597_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s597_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s597_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s597_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s597_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s598_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s598_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s598_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s598_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s598_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s598_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s599_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s599_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s599_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s599_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s599_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s599_val_n5;
    (* src = "src/sreg.spade:138,5" *)
    reg \s600_val ;
    (* src = "src/sreg.spade:138,5" *)
    reg s600_val_n1;
    (* src = "src/sreg.spade:138,5" *)
    reg s600_val_n2;
    (* src = "src/sreg.spade:138,5" *)
    reg s600_val_n3;
    (* src = "src/sreg.spade:138,5" *)
    reg s600_val_n4;
    (* src = "src/sreg.spade:138,5" *)
    reg s600_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg \s601_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s601_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s601_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s601_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s601_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s601_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s601_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s602_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s602_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s602_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s602_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s602_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s602_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s602_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s603_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s603_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s603_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s603_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s603_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s603_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s603_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s604_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s604_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s604_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s604_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s604_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s604_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s604_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s605_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s605_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s605_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s605_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s605_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s605_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s605_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s606_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s606_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s606_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s606_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s606_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s606_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s606_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s607_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s607_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s607_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s607_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s607_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s607_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s607_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s608_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s608_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s608_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s608_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s608_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s608_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s608_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s609_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s609_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s609_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s609_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s609_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s609_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s609_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s610_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s610_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s610_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s610_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s610_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s610_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s610_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s611_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s611_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s611_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s611_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s611_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s611_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s611_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s612_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s612_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s612_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s612_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s612_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s612_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s612_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s613_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s613_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s613_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s613_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s613_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s613_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s613_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s614_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s614_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s614_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s614_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s614_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s614_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s614_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s615_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s615_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s615_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s615_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s615_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s615_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s615_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s616_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s616_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s616_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s616_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s616_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s616_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s616_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s617_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s617_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s617_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s617_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s617_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s617_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s617_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s618_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s618_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s618_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s618_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s618_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s618_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s618_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s619_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s619_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s619_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s619_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s619_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s619_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s619_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s620_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s620_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s620_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s620_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s620_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s620_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s620_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s621_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s621_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s621_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s621_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s621_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s621_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s621_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s622_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s622_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s622_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s622_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s622_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s622_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s622_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s623_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s623_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s623_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s623_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s623_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s623_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s623_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s624_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s624_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s624_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s624_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s624_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s624_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s624_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s625_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s625_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s625_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s625_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s625_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s625_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s625_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s626_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s626_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s626_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s626_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s626_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s626_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s626_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s627_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s627_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s627_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s627_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s627_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s627_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s627_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s628_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s628_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s628_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s628_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s628_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s628_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s628_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s629_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s629_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s629_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s629_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s629_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s629_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s629_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s630_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s630_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s630_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s630_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s630_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s630_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s630_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s631_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s631_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s631_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s631_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s631_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s631_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s631_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s632_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s632_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s632_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s632_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s632_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s632_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s632_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s633_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s633_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s633_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s633_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s633_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s633_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s633_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s634_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s634_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s634_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s634_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s634_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s634_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s634_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s635_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s635_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s635_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s635_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s635_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s635_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s635_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s636_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s636_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s636_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s636_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s636_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s636_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s636_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s637_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s637_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s637_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s637_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s637_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s637_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s637_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s638_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s638_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s638_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s638_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s638_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s638_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s638_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s639_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s639_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s639_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s639_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s639_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s639_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s639_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s640_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s640_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s640_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s640_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s640_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s640_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s640_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s641_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s641_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s641_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s641_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s641_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s641_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s641_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s642_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s642_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s642_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s642_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s642_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s642_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s642_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s643_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s643_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s643_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s643_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s643_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s643_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s643_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s644_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s644_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s644_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s644_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s644_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s644_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s644_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s645_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s645_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s645_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s645_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s645_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s645_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s645_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s646_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s646_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s646_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s646_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s646_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s646_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s646_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s647_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s647_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s647_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s647_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s647_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s647_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s647_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s648_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s648_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s648_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s648_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s648_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s648_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s648_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s649_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s649_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s649_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s649_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s649_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s649_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s649_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s650_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s650_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s650_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s650_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s650_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s650_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s650_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s651_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s651_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s651_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s651_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s651_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s651_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s651_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s652_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s652_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s652_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s652_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s652_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s652_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s652_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s653_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s653_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s653_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s653_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s653_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s653_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s653_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s654_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s654_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s654_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s654_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s654_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s654_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s654_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s655_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s655_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s655_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s655_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s655_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s655_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s655_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s656_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s656_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s656_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s656_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s656_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s656_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s656_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s657_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s657_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s657_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s657_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s657_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s657_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s657_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s658_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s658_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s658_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s658_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s658_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s658_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s658_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s659_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s659_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s659_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s659_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s659_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s659_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s659_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s660_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s660_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s660_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s660_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s660_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s660_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s660_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s661_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s661_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s661_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s661_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s661_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s661_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s661_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s662_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s662_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s662_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s662_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s662_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s662_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s662_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s663_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s663_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s663_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s663_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s663_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s663_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s663_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s664_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s664_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s664_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s664_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s664_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s664_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s664_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s665_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s665_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s665_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s665_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s665_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s665_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s665_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s666_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s666_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s666_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s666_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s666_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s666_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s666_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s667_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s667_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s667_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s667_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s667_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s667_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s667_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s668_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s668_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s668_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s668_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s668_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s668_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s668_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s669_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s669_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s669_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s669_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s669_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s669_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s669_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s670_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s670_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s670_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s670_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s670_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s670_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s670_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s671_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s671_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s671_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s671_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s671_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s671_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s671_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s672_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s672_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s672_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s672_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s672_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s672_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s672_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s673_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s673_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s673_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s673_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s673_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s673_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s673_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s674_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s674_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s674_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s674_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s674_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s674_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s674_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s675_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s675_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s675_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s675_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s675_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s675_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s675_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s676_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s676_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s676_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s676_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s676_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s676_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s676_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s677_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s677_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s677_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s677_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s677_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s677_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s677_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s678_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s678_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s678_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s678_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s678_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s678_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s678_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s679_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s679_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s679_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s679_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s679_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s679_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s679_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s680_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s680_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s680_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s680_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s680_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s680_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s680_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s681_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s681_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s681_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s681_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s681_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s681_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s681_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s682_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s682_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s682_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s682_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s682_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s682_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s682_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s683_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s683_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s683_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s683_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s683_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s683_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s683_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s684_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s684_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s684_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s684_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s684_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s684_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s684_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s685_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s685_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s685_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s685_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s685_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s685_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s685_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s686_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s686_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s686_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s686_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s686_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s686_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s686_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s687_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s687_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s687_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s687_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s687_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s687_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s687_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s688_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s688_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s688_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s688_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s688_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s688_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s688_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s689_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s689_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s689_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s689_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s689_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s689_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s689_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s690_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s690_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s690_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s690_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s690_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s690_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s690_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s691_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s691_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s691_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s691_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s691_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s691_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s691_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s692_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s692_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s692_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s692_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s692_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s692_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s692_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s693_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s693_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s693_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s693_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s693_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s693_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s693_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s694_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s694_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s694_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s694_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s694_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s694_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s694_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s695_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s695_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s695_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s695_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s695_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s695_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s695_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s696_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s696_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s696_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s696_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s696_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s696_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s696_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s697_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s697_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s697_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s697_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s697_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s697_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s697_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s698_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s698_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s698_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s698_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s698_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s698_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s698_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s699_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s699_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s699_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s699_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s699_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s699_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s699_val_n6;
    (* src = "src/sreg.spade:140,5" *)
    reg \s700_val ;
    (* src = "src/sreg.spade:140,5" *)
    reg s700_val_n1;
    (* src = "src/sreg.spade:140,5" *)
    reg s700_val_n2;
    (* src = "src/sreg.spade:140,5" *)
    reg s700_val_n3;
    (* src = "src/sreg.spade:140,5" *)
    reg s700_val_n4;
    (* src = "src/sreg.spade:140,5" *)
    reg s700_val_n5;
    (* src = "src/sreg.spade:140,5" *)
    reg s700_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg \s701_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s701_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s701_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s701_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s701_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s701_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s701_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s701_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s702_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s702_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s702_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s702_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s702_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s702_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s702_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s702_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s703_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s703_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s703_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s703_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s703_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s703_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s703_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s703_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s704_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s704_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s704_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s704_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s704_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s704_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s704_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s704_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s705_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s705_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s705_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s705_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s705_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s705_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s705_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s705_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s706_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s706_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s706_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s706_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s706_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s706_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s706_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s706_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s707_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s707_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s707_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s707_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s707_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s707_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s707_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s707_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s708_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s708_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s708_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s708_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s708_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s708_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s708_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s708_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s709_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s709_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s709_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s709_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s709_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s709_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s709_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s709_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s710_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s710_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s710_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s710_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s710_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s710_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s710_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s710_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s711_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s711_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s711_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s711_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s711_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s711_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s711_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s711_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s712_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s712_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s712_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s712_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s712_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s712_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s712_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s712_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s713_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s713_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s713_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s713_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s713_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s713_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s713_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s713_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s714_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s714_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s714_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s714_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s714_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s714_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s714_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s714_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s715_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s715_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s715_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s715_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s715_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s715_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s715_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s715_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s716_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s716_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s716_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s716_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s716_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s716_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s716_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s716_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s717_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s717_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s717_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s717_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s717_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s717_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s717_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s717_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s718_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s718_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s718_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s718_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s718_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s718_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s718_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s718_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s719_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s719_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s719_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s719_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s719_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s719_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s719_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s719_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s720_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s720_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s720_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s720_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s720_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s720_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s720_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s720_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s721_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s721_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s721_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s721_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s721_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s721_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s721_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s721_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s722_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s722_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s722_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s722_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s722_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s722_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s722_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s722_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s723_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s723_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s723_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s723_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s723_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s723_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s723_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s723_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s724_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s724_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s724_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s724_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s724_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s724_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s724_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s724_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s725_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s725_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s725_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s725_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s725_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s725_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s725_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s725_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s726_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s726_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s726_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s726_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s726_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s726_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s726_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s726_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s727_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s727_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s727_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s727_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s727_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s727_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s727_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s727_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s728_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s728_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s728_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s728_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s728_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s728_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s728_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s728_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s729_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s729_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s729_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s729_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s729_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s729_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s729_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s729_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s730_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s730_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s730_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s730_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s730_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s730_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s730_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s730_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s731_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s731_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s731_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s731_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s731_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s731_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s731_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s731_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s732_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s732_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s732_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s732_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s732_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s732_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s732_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s732_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s733_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s733_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s733_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s733_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s733_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s733_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s733_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s733_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s734_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s734_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s734_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s734_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s734_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s734_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s734_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s734_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s735_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s735_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s735_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s735_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s735_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s735_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s735_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s735_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s736_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s736_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s736_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s736_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s736_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s736_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s736_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s736_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s737_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s737_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s737_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s737_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s737_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s737_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s737_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s737_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s738_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s738_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s738_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s738_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s738_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s738_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s738_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s738_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s739_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s739_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s739_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s739_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s739_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s739_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s739_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s739_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s740_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s740_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s740_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s740_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s740_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s740_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s740_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s740_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s741_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s741_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s741_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s741_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s741_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s741_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s741_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s741_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s742_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s742_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s742_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s742_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s742_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s742_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s742_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s742_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s743_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s743_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s743_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s743_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s743_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s743_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s743_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s743_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s744_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s744_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s744_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s744_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s744_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s744_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s744_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s744_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s745_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s745_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s745_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s745_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s745_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s745_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s745_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s745_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s746_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s746_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s746_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s746_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s746_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s746_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s746_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s746_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s747_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s747_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s747_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s747_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s747_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s747_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s747_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s747_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s748_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s748_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s748_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s748_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s748_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s748_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s748_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s748_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s749_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s749_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s749_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s749_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s749_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s749_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s749_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s749_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s750_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s750_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s750_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s750_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s750_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s750_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s750_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s750_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s751_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s751_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s751_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s751_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s751_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s751_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s751_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s751_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s752_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s752_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s752_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s752_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s752_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s752_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s752_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s752_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s753_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s753_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s753_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s753_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s753_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s753_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s753_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s753_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s754_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s754_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s754_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s754_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s754_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s754_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s754_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s754_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s755_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s755_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s755_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s755_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s755_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s755_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s755_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s755_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s756_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s756_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s756_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s756_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s756_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s756_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s756_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s756_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s757_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s757_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s757_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s757_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s757_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s757_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s757_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s757_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s758_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s758_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s758_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s758_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s758_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s758_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s758_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s758_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s759_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s759_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s759_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s759_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s759_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s759_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s759_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s759_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s760_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s760_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s760_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s760_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s760_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s760_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s760_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s760_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s761_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s761_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s761_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s761_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s761_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s761_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s761_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s761_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s762_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s762_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s762_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s762_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s762_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s762_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s762_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s762_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s763_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s763_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s763_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s763_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s763_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s763_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s763_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s763_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s764_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s764_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s764_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s764_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s764_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s764_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s764_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s764_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s765_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s765_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s765_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s765_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s765_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s765_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s765_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s765_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s766_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s766_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s766_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s766_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s766_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s766_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s766_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s766_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s767_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s767_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s767_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s767_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s767_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s767_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s767_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s767_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s768_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s768_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s768_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s768_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s768_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s768_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s768_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s768_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s769_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s769_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s769_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s769_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s769_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s769_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s769_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s769_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s770_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s770_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s770_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s770_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s770_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s770_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s770_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s770_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s771_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s771_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s771_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s771_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s771_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s771_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s771_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s771_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s772_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s772_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s772_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s772_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s772_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s772_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s772_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s772_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s773_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s773_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s773_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s773_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s773_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s773_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s773_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s773_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s774_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s774_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s774_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s774_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s774_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s774_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s774_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s774_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s775_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s775_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s775_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s775_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s775_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s775_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s775_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s775_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s776_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s776_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s776_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s776_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s776_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s776_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s776_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s776_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s777_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s777_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s777_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s777_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s777_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s777_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s777_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s777_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s778_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s778_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s778_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s778_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s778_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s778_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s778_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s778_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s779_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s779_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s779_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s779_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s779_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s779_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s779_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s779_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s780_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s780_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s780_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s780_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s780_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s780_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s780_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s780_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s781_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s781_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s781_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s781_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s781_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s781_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s781_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s781_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s782_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s782_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s782_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s782_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s782_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s782_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s782_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s782_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s783_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s783_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s783_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s783_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s783_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s783_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s783_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s783_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s784_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s784_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s784_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s784_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s784_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s784_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s784_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s784_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s785_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s785_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s785_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s785_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s785_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s785_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s785_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s785_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s786_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s786_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s786_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s786_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s786_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s786_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s786_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s786_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s787_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s787_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s787_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s787_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s787_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s787_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s787_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s787_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s788_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s788_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s788_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s788_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s788_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s788_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s788_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s788_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s789_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s789_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s789_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s789_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s789_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s789_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s789_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s789_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s790_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s790_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s790_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s790_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s790_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s790_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s790_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s790_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s791_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s791_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s791_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s791_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s791_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s791_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s791_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s791_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s792_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s792_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s792_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s792_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s792_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s792_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s792_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s792_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s793_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s793_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s793_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s793_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s793_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s793_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s793_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s793_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s794_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s794_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s794_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s794_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s794_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s794_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s794_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s794_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s795_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s795_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s795_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s795_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s795_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s795_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s795_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s795_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s796_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s796_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s796_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s796_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s796_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s796_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s796_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s796_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s797_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s797_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s797_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s797_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s797_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s797_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s797_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s797_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s798_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s798_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s798_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s798_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s798_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s798_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s798_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s798_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s799_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s799_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s799_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s799_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s799_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s799_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s799_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s799_val_n7;
    (* src = "src/sreg.spade:142,5" *)
    reg \s800_val ;
    (* src = "src/sreg.spade:142,5" *)
    reg s800_val_n1;
    (* src = "src/sreg.spade:142,5" *)
    reg s800_val_n2;
    (* src = "src/sreg.spade:142,5" *)
    reg s800_val_n3;
    (* src = "src/sreg.spade:142,5" *)
    reg s800_val_n4;
    (* src = "src/sreg.spade:142,5" *)
    reg s800_val_n5;
    (* src = "src/sreg.spade:142,5" *)
    reg s800_val_n6;
    (* src = "src/sreg.spade:142,5" *)
    reg s800_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg \s801_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s801_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s801_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s801_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s801_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s801_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s801_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s801_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s801_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s802_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s802_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s802_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s802_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s802_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s802_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s802_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s802_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s802_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s803_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s803_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s803_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s803_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s803_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s803_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s803_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s803_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s803_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s804_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s804_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s804_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s804_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s804_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s804_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s804_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s804_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s804_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s805_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s805_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s805_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s805_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s805_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s805_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s805_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s805_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s805_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s806_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s806_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s806_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s806_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s806_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s806_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s806_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s806_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s806_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s807_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s807_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s807_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s807_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s807_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s807_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s807_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s807_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s807_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s808_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s808_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s808_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s808_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s808_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s808_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s808_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s808_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s808_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s809_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s809_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s809_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s809_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s809_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s809_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s809_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s809_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s809_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s810_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s810_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s810_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s810_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s810_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s810_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s810_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s810_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s810_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s811_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s811_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s811_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s811_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s811_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s811_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s811_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s811_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s811_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s812_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s812_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s812_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s812_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s812_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s812_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s812_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s812_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s812_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s813_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s813_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s813_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s813_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s813_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s813_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s813_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s813_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s813_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s814_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s814_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s814_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s814_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s814_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s814_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s814_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s814_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s814_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s815_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s815_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s815_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s815_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s815_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s815_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s815_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s815_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s815_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s816_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s816_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s816_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s816_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s816_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s816_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s816_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s816_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s816_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s817_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s817_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s817_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s817_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s817_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s817_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s817_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s817_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s817_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s818_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s818_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s818_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s818_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s818_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s818_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s818_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s818_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s818_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s819_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s819_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s819_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s819_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s819_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s819_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s819_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s819_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s819_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s820_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s820_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s820_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s820_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s820_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s820_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s820_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s820_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s820_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s821_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s821_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s821_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s821_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s821_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s821_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s821_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s821_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s821_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s822_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s822_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s822_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s822_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s822_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s822_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s822_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s822_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s822_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s823_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s823_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s823_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s823_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s823_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s823_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s823_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s823_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s823_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s824_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s824_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s824_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s824_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s824_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s824_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s824_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s824_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s824_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s825_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s825_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s825_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s825_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s825_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s825_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s825_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s825_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s825_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s826_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s826_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s826_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s826_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s826_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s826_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s826_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s826_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s826_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s827_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s827_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s827_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s827_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s827_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s827_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s827_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s827_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s827_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s828_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s828_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s828_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s828_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s828_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s828_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s828_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s828_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s828_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s829_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s829_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s829_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s829_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s829_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s829_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s829_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s829_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s829_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s830_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s830_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s830_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s830_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s830_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s830_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s830_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s830_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s830_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s831_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s831_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s831_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s831_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s831_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s831_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s831_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s831_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s831_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s832_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s832_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s832_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s832_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s832_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s832_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s832_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s832_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s832_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s833_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s833_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s833_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s833_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s833_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s833_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s833_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s833_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s833_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s834_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s834_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s834_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s834_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s834_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s834_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s834_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s834_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s834_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s835_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s835_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s835_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s835_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s835_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s835_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s835_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s835_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s835_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s836_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s836_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s836_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s836_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s836_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s836_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s836_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s836_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s836_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s837_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s837_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s837_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s837_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s837_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s837_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s837_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s837_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s837_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s838_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s838_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s838_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s838_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s838_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s838_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s838_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s838_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s838_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s839_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s839_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s839_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s839_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s839_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s839_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s839_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s839_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s839_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s840_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s840_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s840_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s840_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s840_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s840_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s840_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s840_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s840_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s841_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s841_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s841_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s841_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s841_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s841_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s841_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s841_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s841_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s842_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s842_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s842_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s842_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s842_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s842_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s842_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s842_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s842_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s843_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s843_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s843_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s843_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s843_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s843_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s843_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s843_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s843_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s844_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s844_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s844_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s844_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s844_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s844_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s844_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s844_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s844_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s845_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s845_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s845_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s845_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s845_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s845_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s845_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s845_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s845_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s846_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s846_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s846_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s846_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s846_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s846_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s846_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s846_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s846_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s847_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s847_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s847_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s847_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s847_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s847_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s847_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s847_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s847_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s848_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s848_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s848_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s848_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s848_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s848_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s848_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s848_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s848_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s849_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s849_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s849_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s849_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s849_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s849_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s849_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s849_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s849_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s850_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s850_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s850_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s850_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s850_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s850_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s850_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s850_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s850_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s851_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s851_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s851_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s851_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s851_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s851_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s851_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s851_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s851_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s852_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s852_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s852_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s852_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s852_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s852_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s852_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s852_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s852_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s853_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s853_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s853_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s853_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s853_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s853_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s853_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s853_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s853_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s854_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s854_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s854_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s854_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s854_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s854_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s854_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s854_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s854_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s855_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s855_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s855_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s855_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s855_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s855_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s855_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s855_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s855_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s856_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s856_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s856_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s856_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s856_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s856_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s856_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s856_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s856_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s857_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s857_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s857_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s857_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s857_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s857_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s857_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s857_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s857_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s858_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s858_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s858_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s858_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s858_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s858_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s858_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s858_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s858_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s859_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s859_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s859_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s859_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s859_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s859_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s859_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s859_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s859_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s860_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s860_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s860_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s860_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s860_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s860_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s860_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s860_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s860_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s861_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s861_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s861_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s861_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s861_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s861_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s861_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s861_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s861_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s862_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s862_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s862_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s862_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s862_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s862_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s862_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s862_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s862_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s863_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s863_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s863_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s863_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s863_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s863_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s863_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s863_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s863_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s864_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s864_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s864_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s864_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s864_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s864_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s864_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s864_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s864_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s865_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s865_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s865_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s865_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s865_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s865_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s865_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s865_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s865_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s866_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s866_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s866_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s866_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s866_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s866_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s866_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s866_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s866_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s867_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s867_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s867_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s867_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s867_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s867_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s867_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s867_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s867_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s868_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s868_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s868_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s868_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s868_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s868_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s868_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s868_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s868_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s869_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s869_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s869_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s869_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s869_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s869_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s869_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s869_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s869_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s870_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s870_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s870_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s870_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s870_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s870_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s870_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s870_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s870_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s871_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s871_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s871_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s871_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s871_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s871_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s871_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s871_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s871_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s872_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s872_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s872_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s872_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s872_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s872_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s872_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s872_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s872_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s873_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s873_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s873_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s873_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s873_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s873_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s873_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s873_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s873_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s874_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s874_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s874_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s874_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s874_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s874_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s874_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s874_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s874_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s875_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s875_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s875_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s875_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s875_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s875_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s875_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s875_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s875_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s876_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s876_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s876_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s876_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s876_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s876_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s876_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s876_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s876_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s877_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s877_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s877_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s877_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s877_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s877_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s877_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s877_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s877_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s878_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s878_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s878_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s878_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s878_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s878_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s878_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s878_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s878_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s879_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s879_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s879_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s879_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s879_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s879_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s879_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s879_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s879_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s880_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s880_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s880_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s880_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s880_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s880_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s880_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s880_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s880_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s881_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s881_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s881_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s881_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s881_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s881_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s881_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s881_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s881_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s882_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s882_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s882_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s882_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s882_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s882_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s882_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s882_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s882_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s883_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s883_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s883_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s883_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s883_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s883_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s883_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s883_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s883_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s884_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s884_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s884_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s884_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s884_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s884_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s884_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s884_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s884_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s885_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s885_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s885_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s885_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s885_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s885_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s885_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s885_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s885_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s886_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s886_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s886_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s886_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s886_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s886_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s886_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s886_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s886_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s887_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s887_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s887_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s887_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s887_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s887_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s887_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s887_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s887_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s888_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s888_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s888_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s888_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s888_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s888_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s888_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s888_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s888_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s889_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s889_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s889_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s889_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s889_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s889_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s889_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s889_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s889_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s890_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s890_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s890_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s890_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s890_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s890_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s890_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s890_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s890_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s891_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s891_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s891_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s891_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s891_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s891_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s891_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s891_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s891_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s892_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s892_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s892_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s892_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s892_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s892_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s892_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s892_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s892_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s893_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s893_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s893_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s893_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s893_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s893_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s893_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s893_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s893_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s894_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s894_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s894_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s894_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s894_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s894_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s894_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s894_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s894_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s895_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s895_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s895_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s895_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s895_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s895_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s895_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s895_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s895_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s896_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s896_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s896_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s896_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s896_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s896_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s896_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s896_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s896_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s897_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s897_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s897_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s897_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s897_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s897_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s897_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s897_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s897_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s898_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s898_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s898_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s898_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s898_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s898_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s898_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s898_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s898_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s899_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s899_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s899_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s899_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s899_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s899_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s899_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s899_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s899_val_n8;
    (* src = "src/sreg.spade:144,5" *)
    reg \s900_val ;
    (* src = "src/sreg.spade:144,5" *)
    reg s900_val_n1;
    (* src = "src/sreg.spade:144,5" *)
    reg s900_val_n2;
    (* src = "src/sreg.spade:144,5" *)
    reg s900_val_n3;
    (* src = "src/sreg.spade:144,5" *)
    reg s900_val_n4;
    (* src = "src/sreg.spade:144,5" *)
    reg s900_val_n5;
    (* src = "src/sreg.spade:144,5" *)
    reg s900_val_n6;
    (* src = "src/sreg.spade:144,5" *)
    reg s900_val_n7;
    (* src = "src/sreg.spade:144,5" *)
    reg s900_val_n8;
    (* src = "src/sreg.spade:127,19" *)
    logic val_n1;
    (* src = "src/sreg.spade:129,19" *)
    logic val_n2;
    (* src = "src/sreg.spade:131,19" *)
    logic val_n3;
    (* src = "src/sreg.spade:133,19" *)
    logic val_n4;
    (* src = "src/sreg.spade:135,19" *)
    logic val_n5;
    (* src = "src/sreg.spade:137,19" *)
    logic val_n6;
    (* src = "src/sreg.spade:139,19" *)
    logic val_n7;
    (* src = "src/sreg.spade:141,19" *)
    logic val_n8;
    (* src = "src/sreg.spade:143,19" *)
    logic val_n9;
    always @(posedge \clk ) begin
        \s1_val  <= \val ;
    end
    always @(posedge \clk ) begin
        \s2_val  <= \s1_val ;
    end
    always @(posedge \clk ) begin
        \s3_val  <= \s2_val ;
    end
    always @(posedge \clk ) begin
        \s4_val  <= \s3_val ;
    end
    always @(posedge \clk ) begin
        \s5_val  <= \s4_val ;
    end
    always @(posedge \clk ) begin
        \s6_val  <= \s5_val ;
    end
    always @(posedge \clk ) begin
        \s7_val  <= \s6_val ;
    end
    always @(posedge \clk ) begin
        \s8_val  <= \s7_val ;
    end
    always @(posedge \clk ) begin
        \s9_val  <= \s8_val ;
    end
    always @(posedge \clk ) begin
        \s10_val  <= \s9_val ;
    end
    always @(posedge \clk ) begin
        \s11_val  <= \s10_val ;
    end
    always @(posedge \clk ) begin
        \s12_val  <= \s11_val ;
    end
    always @(posedge \clk ) begin
        \s13_val  <= \s12_val ;
    end
    always @(posedge \clk ) begin
        \s14_val  <= \s13_val ;
    end
    always @(posedge \clk ) begin
        \s15_val  <= \s14_val ;
    end
    always @(posedge \clk ) begin
        \s16_val  <= \s15_val ;
    end
    always @(posedge \clk ) begin
        \s17_val  <= \s16_val ;
    end
    always @(posedge \clk ) begin
        \s18_val  <= \s17_val ;
    end
    always @(posedge \clk ) begin
        \s19_val  <= \s18_val ;
    end
    always @(posedge \clk ) begin
        \s20_val  <= \s19_val ;
    end
    always @(posedge \clk ) begin
        \s21_val  <= \s20_val ;
    end
    always @(posedge \clk ) begin
        \s22_val  <= \s21_val ;
    end
    always @(posedge \clk ) begin
        \s23_val  <= \s22_val ;
    end
    always @(posedge \clk ) begin
        \s24_val  <= \s23_val ;
    end
    always @(posedge \clk ) begin
        \s25_val  <= \s24_val ;
    end
    always @(posedge \clk ) begin
        \s26_val  <= \s25_val ;
    end
    always @(posedge \clk ) begin
        \s27_val  <= \s26_val ;
    end
    always @(posedge \clk ) begin
        \s28_val  <= \s27_val ;
    end
    always @(posedge \clk ) begin
        \s29_val  <= \s28_val ;
    end
    always @(posedge \clk ) begin
        \s30_val  <= \s29_val ;
    end
    always @(posedge \clk ) begin
        \s31_val  <= \s30_val ;
    end
    always @(posedge \clk ) begin
        \s32_val  <= \s31_val ;
    end
    always @(posedge \clk ) begin
        \s33_val  <= \s32_val ;
    end
    always @(posedge \clk ) begin
        \s34_val  <= \s33_val ;
    end
    always @(posedge \clk ) begin
        \s35_val  <= \s34_val ;
    end
    always @(posedge \clk ) begin
        \s36_val  <= \s35_val ;
    end
    always @(posedge \clk ) begin
        \s37_val  <= \s36_val ;
    end
    always @(posedge \clk ) begin
        \s38_val  <= \s37_val ;
    end
    always @(posedge \clk ) begin
        \s39_val  <= \s38_val ;
    end
    always @(posedge \clk ) begin
        \s40_val  <= \s39_val ;
    end
    always @(posedge \clk ) begin
        \s41_val  <= \s40_val ;
    end
    always @(posedge \clk ) begin
        \s42_val  <= \s41_val ;
    end
    always @(posedge \clk ) begin
        \s43_val  <= \s42_val ;
    end
    always @(posedge \clk ) begin
        \s44_val  <= \s43_val ;
    end
    always @(posedge \clk ) begin
        \s45_val  <= \s44_val ;
    end
    always @(posedge \clk ) begin
        \s46_val  <= \s45_val ;
    end
    always @(posedge \clk ) begin
        \s47_val  <= \s46_val ;
    end
    always @(posedge \clk ) begin
        \s48_val  <= \s47_val ;
    end
    always @(posedge \clk ) begin
        \s49_val  <= \s48_val ;
    end
    always @(posedge \clk ) begin
        \s50_val  <= \s49_val ;
    end
    always @(posedge \clk ) begin
        \s51_val  <= \s50_val ;
    end
    always @(posedge \clk ) begin
        \s52_val  <= \s51_val ;
    end
    always @(posedge \clk ) begin
        \s53_val  <= \s52_val ;
    end
    always @(posedge \clk ) begin
        \s54_val  <= \s53_val ;
    end
    always @(posedge \clk ) begin
        \s55_val  <= \s54_val ;
    end
    always @(posedge \clk ) begin
        \s56_val  <= \s55_val ;
    end
    always @(posedge \clk ) begin
        \s57_val  <= \s56_val ;
    end
    always @(posedge \clk ) begin
        \s58_val  <= \s57_val ;
    end
    always @(posedge \clk ) begin
        \s59_val  <= \s58_val ;
    end
    always @(posedge \clk ) begin
        \s60_val  <= \s59_val ;
    end
    always @(posedge \clk ) begin
        \s61_val  <= \s60_val ;
    end
    always @(posedge \clk ) begin
        \s62_val  <= \s61_val ;
    end
    always @(posedge \clk ) begin
        \s63_val  <= \s62_val ;
    end
    always @(posedge \clk ) begin
        \s64_val  <= \s63_val ;
    end
    always @(posedge \clk ) begin
        \s65_val  <= \s64_val ;
    end
    always @(posedge \clk ) begin
        \s66_val  <= \s65_val ;
    end
    always @(posedge \clk ) begin
        \s67_val  <= \s66_val ;
    end
    always @(posedge \clk ) begin
        \s68_val  <= \s67_val ;
    end
    always @(posedge \clk ) begin
        \s69_val  <= \s68_val ;
    end
    always @(posedge \clk ) begin
        \s70_val  <= \s69_val ;
    end
    always @(posedge \clk ) begin
        \s71_val  <= \s70_val ;
    end
    always @(posedge \clk ) begin
        \s72_val  <= \s71_val ;
    end
    always @(posedge \clk ) begin
        \s73_val  <= \s72_val ;
    end
    always @(posedge \clk ) begin
        \s74_val  <= \s73_val ;
    end
    always @(posedge \clk ) begin
        \s75_val  <= \s74_val ;
    end
    always @(posedge \clk ) begin
        \s76_val  <= \s75_val ;
    end
    always @(posedge \clk ) begin
        \s77_val  <= \s76_val ;
    end
    always @(posedge \clk ) begin
        \s78_val  <= \s77_val ;
    end
    always @(posedge \clk ) begin
        \s79_val  <= \s78_val ;
    end
    always @(posedge \clk ) begin
        \s80_val  <= \s79_val ;
    end
    always @(posedge \clk ) begin
        \s81_val  <= \s80_val ;
    end
    always @(posedge \clk ) begin
        \s82_val  <= \s81_val ;
    end
    always @(posedge \clk ) begin
        \s83_val  <= \s82_val ;
    end
    always @(posedge \clk ) begin
        \s84_val  <= \s83_val ;
    end
    always @(posedge \clk ) begin
        \s85_val  <= \s84_val ;
    end
    always @(posedge \clk ) begin
        \s86_val  <= \s85_val ;
    end
    always @(posedge \clk ) begin
        \s87_val  <= \s86_val ;
    end
    always @(posedge \clk ) begin
        \s88_val  <= \s87_val ;
    end
    always @(posedge \clk ) begin
        \s89_val  <= \s88_val ;
    end
    always @(posedge \clk ) begin
        \s90_val  <= \s89_val ;
    end
    always @(posedge \clk ) begin
        \s91_val  <= \s90_val ;
    end
    always @(posedge \clk ) begin
        \s92_val  <= \s91_val ;
    end
    always @(posedge \clk ) begin
        \s93_val  <= \s92_val ;
    end
    always @(posedge \clk ) begin
        \s94_val  <= \s93_val ;
    end
    always @(posedge \clk ) begin
        \s95_val  <= \s94_val ;
    end
    always @(posedge \clk ) begin
        \s96_val  <= \s95_val ;
    end
    always @(posedge \clk ) begin
        \s97_val  <= \s96_val ;
    end
    always @(posedge \clk ) begin
        \s98_val  <= \s97_val ;
    end
    always @(posedge \clk ) begin
        \s99_val  <= \s98_val ;
    end
    always @(posedge \clk ) begin
        \s100_val  <= \s99_val ;
    end
    always @(posedge \clk ) begin
        \s101_val  <= \s100_val ;
    end
    always @(posedge \clk ) begin
        s101_val_n1 <= val_n1;
    end
    always @(posedge \clk ) begin
        \s102_val  <= \s101_val ;
    end
    always @(posedge \clk ) begin
        s102_val_n1 <= s101_val_n1;
    end
    always @(posedge \clk ) begin
        \s103_val  <= \s102_val ;
    end
    always @(posedge \clk ) begin
        s103_val_n1 <= s102_val_n1;
    end
    always @(posedge \clk ) begin
        \s104_val  <= \s103_val ;
    end
    always @(posedge \clk ) begin
        s104_val_n1 <= s103_val_n1;
    end
    always @(posedge \clk ) begin
        \s105_val  <= \s104_val ;
    end
    always @(posedge \clk ) begin
        s105_val_n1 <= s104_val_n1;
    end
    always @(posedge \clk ) begin
        \s106_val  <= \s105_val ;
    end
    always @(posedge \clk ) begin
        s106_val_n1 <= s105_val_n1;
    end
    always @(posedge \clk ) begin
        \s107_val  <= \s106_val ;
    end
    always @(posedge \clk ) begin
        s107_val_n1 <= s106_val_n1;
    end
    always @(posedge \clk ) begin
        \s108_val  <= \s107_val ;
    end
    always @(posedge \clk ) begin
        s108_val_n1 <= s107_val_n1;
    end
    always @(posedge \clk ) begin
        \s109_val  <= \s108_val ;
    end
    always @(posedge \clk ) begin
        s109_val_n1 <= s108_val_n1;
    end
    always @(posedge \clk ) begin
        \s110_val  <= \s109_val ;
    end
    always @(posedge \clk ) begin
        s110_val_n1 <= s109_val_n1;
    end
    always @(posedge \clk ) begin
        \s111_val  <= \s110_val ;
    end
    always @(posedge \clk ) begin
        s111_val_n1 <= s110_val_n1;
    end
    always @(posedge \clk ) begin
        \s112_val  <= \s111_val ;
    end
    always @(posedge \clk ) begin
        s112_val_n1 <= s111_val_n1;
    end
    always @(posedge \clk ) begin
        \s113_val  <= \s112_val ;
    end
    always @(posedge \clk ) begin
        s113_val_n1 <= s112_val_n1;
    end
    always @(posedge \clk ) begin
        \s114_val  <= \s113_val ;
    end
    always @(posedge \clk ) begin
        s114_val_n1 <= s113_val_n1;
    end
    always @(posedge \clk ) begin
        \s115_val  <= \s114_val ;
    end
    always @(posedge \clk ) begin
        s115_val_n1 <= s114_val_n1;
    end
    always @(posedge \clk ) begin
        \s116_val  <= \s115_val ;
    end
    always @(posedge \clk ) begin
        s116_val_n1 <= s115_val_n1;
    end
    always @(posedge \clk ) begin
        \s117_val  <= \s116_val ;
    end
    always @(posedge \clk ) begin
        s117_val_n1 <= s116_val_n1;
    end
    always @(posedge \clk ) begin
        \s118_val  <= \s117_val ;
    end
    always @(posedge \clk ) begin
        s118_val_n1 <= s117_val_n1;
    end
    always @(posedge \clk ) begin
        \s119_val  <= \s118_val ;
    end
    always @(posedge \clk ) begin
        s119_val_n1 <= s118_val_n1;
    end
    always @(posedge \clk ) begin
        \s120_val  <= \s119_val ;
    end
    always @(posedge \clk ) begin
        s120_val_n1 <= s119_val_n1;
    end
    always @(posedge \clk ) begin
        \s121_val  <= \s120_val ;
    end
    always @(posedge \clk ) begin
        s121_val_n1 <= s120_val_n1;
    end
    always @(posedge \clk ) begin
        \s122_val  <= \s121_val ;
    end
    always @(posedge \clk ) begin
        s122_val_n1 <= s121_val_n1;
    end
    always @(posedge \clk ) begin
        \s123_val  <= \s122_val ;
    end
    always @(posedge \clk ) begin
        s123_val_n1 <= s122_val_n1;
    end
    always @(posedge \clk ) begin
        \s124_val  <= \s123_val ;
    end
    always @(posedge \clk ) begin
        s124_val_n1 <= s123_val_n1;
    end
    always @(posedge \clk ) begin
        \s125_val  <= \s124_val ;
    end
    always @(posedge \clk ) begin
        s125_val_n1 <= s124_val_n1;
    end
    always @(posedge \clk ) begin
        \s126_val  <= \s125_val ;
    end
    always @(posedge \clk ) begin
        s126_val_n1 <= s125_val_n1;
    end
    always @(posedge \clk ) begin
        \s127_val  <= \s126_val ;
    end
    always @(posedge \clk ) begin
        s127_val_n1 <= s126_val_n1;
    end
    always @(posedge \clk ) begin
        \s128_val  <= \s127_val ;
    end
    always @(posedge \clk ) begin
        s128_val_n1 <= s127_val_n1;
    end
    always @(posedge \clk ) begin
        \s129_val  <= \s128_val ;
    end
    always @(posedge \clk ) begin
        s129_val_n1 <= s128_val_n1;
    end
    always @(posedge \clk ) begin
        \s130_val  <= \s129_val ;
    end
    always @(posedge \clk ) begin
        s130_val_n1 <= s129_val_n1;
    end
    always @(posedge \clk ) begin
        \s131_val  <= \s130_val ;
    end
    always @(posedge \clk ) begin
        s131_val_n1 <= s130_val_n1;
    end
    always @(posedge \clk ) begin
        \s132_val  <= \s131_val ;
    end
    always @(posedge \clk ) begin
        s132_val_n1 <= s131_val_n1;
    end
    always @(posedge \clk ) begin
        \s133_val  <= \s132_val ;
    end
    always @(posedge \clk ) begin
        s133_val_n1 <= s132_val_n1;
    end
    always @(posedge \clk ) begin
        \s134_val  <= \s133_val ;
    end
    always @(posedge \clk ) begin
        s134_val_n1 <= s133_val_n1;
    end
    always @(posedge \clk ) begin
        \s135_val  <= \s134_val ;
    end
    always @(posedge \clk ) begin
        s135_val_n1 <= s134_val_n1;
    end
    always @(posedge \clk ) begin
        \s136_val  <= \s135_val ;
    end
    always @(posedge \clk ) begin
        s136_val_n1 <= s135_val_n1;
    end
    always @(posedge \clk ) begin
        \s137_val  <= \s136_val ;
    end
    always @(posedge \clk ) begin
        s137_val_n1 <= s136_val_n1;
    end
    always @(posedge \clk ) begin
        \s138_val  <= \s137_val ;
    end
    always @(posedge \clk ) begin
        s138_val_n1 <= s137_val_n1;
    end
    always @(posedge \clk ) begin
        \s139_val  <= \s138_val ;
    end
    always @(posedge \clk ) begin
        s139_val_n1 <= s138_val_n1;
    end
    always @(posedge \clk ) begin
        \s140_val  <= \s139_val ;
    end
    always @(posedge \clk ) begin
        s140_val_n1 <= s139_val_n1;
    end
    always @(posedge \clk ) begin
        \s141_val  <= \s140_val ;
    end
    always @(posedge \clk ) begin
        s141_val_n1 <= s140_val_n1;
    end
    always @(posedge \clk ) begin
        \s142_val  <= \s141_val ;
    end
    always @(posedge \clk ) begin
        s142_val_n1 <= s141_val_n1;
    end
    always @(posedge \clk ) begin
        \s143_val  <= \s142_val ;
    end
    always @(posedge \clk ) begin
        s143_val_n1 <= s142_val_n1;
    end
    always @(posedge \clk ) begin
        \s144_val  <= \s143_val ;
    end
    always @(posedge \clk ) begin
        s144_val_n1 <= s143_val_n1;
    end
    always @(posedge \clk ) begin
        \s145_val  <= \s144_val ;
    end
    always @(posedge \clk ) begin
        s145_val_n1 <= s144_val_n1;
    end
    always @(posedge \clk ) begin
        \s146_val  <= \s145_val ;
    end
    always @(posedge \clk ) begin
        s146_val_n1 <= s145_val_n1;
    end
    always @(posedge \clk ) begin
        \s147_val  <= \s146_val ;
    end
    always @(posedge \clk ) begin
        s147_val_n1 <= s146_val_n1;
    end
    always @(posedge \clk ) begin
        \s148_val  <= \s147_val ;
    end
    always @(posedge \clk ) begin
        s148_val_n1 <= s147_val_n1;
    end
    always @(posedge \clk ) begin
        \s149_val  <= \s148_val ;
    end
    always @(posedge \clk ) begin
        s149_val_n1 <= s148_val_n1;
    end
    always @(posedge \clk ) begin
        \s150_val  <= \s149_val ;
    end
    always @(posedge \clk ) begin
        s150_val_n1 <= s149_val_n1;
    end
    always @(posedge \clk ) begin
        \s151_val  <= \s150_val ;
    end
    always @(posedge \clk ) begin
        s151_val_n1 <= s150_val_n1;
    end
    always @(posedge \clk ) begin
        \s152_val  <= \s151_val ;
    end
    always @(posedge \clk ) begin
        s152_val_n1 <= s151_val_n1;
    end
    always @(posedge \clk ) begin
        \s153_val  <= \s152_val ;
    end
    always @(posedge \clk ) begin
        s153_val_n1 <= s152_val_n1;
    end
    always @(posedge \clk ) begin
        \s154_val  <= \s153_val ;
    end
    always @(posedge \clk ) begin
        s154_val_n1 <= s153_val_n1;
    end
    always @(posedge \clk ) begin
        \s155_val  <= \s154_val ;
    end
    always @(posedge \clk ) begin
        s155_val_n1 <= s154_val_n1;
    end
    always @(posedge \clk ) begin
        \s156_val  <= \s155_val ;
    end
    always @(posedge \clk ) begin
        s156_val_n1 <= s155_val_n1;
    end
    always @(posedge \clk ) begin
        \s157_val  <= \s156_val ;
    end
    always @(posedge \clk ) begin
        s157_val_n1 <= s156_val_n1;
    end
    always @(posedge \clk ) begin
        \s158_val  <= \s157_val ;
    end
    always @(posedge \clk ) begin
        s158_val_n1 <= s157_val_n1;
    end
    always @(posedge \clk ) begin
        \s159_val  <= \s158_val ;
    end
    always @(posedge \clk ) begin
        s159_val_n1 <= s158_val_n1;
    end
    always @(posedge \clk ) begin
        \s160_val  <= \s159_val ;
    end
    always @(posedge \clk ) begin
        s160_val_n1 <= s159_val_n1;
    end
    always @(posedge \clk ) begin
        \s161_val  <= \s160_val ;
    end
    always @(posedge \clk ) begin
        s161_val_n1 <= s160_val_n1;
    end
    always @(posedge \clk ) begin
        \s162_val  <= \s161_val ;
    end
    always @(posedge \clk ) begin
        s162_val_n1 <= s161_val_n1;
    end
    always @(posedge \clk ) begin
        \s163_val  <= \s162_val ;
    end
    always @(posedge \clk ) begin
        s163_val_n1 <= s162_val_n1;
    end
    always @(posedge \clk ) begin
        \s164_val  <= \s163_val ;
    end
    always @(posedge \clk ) begin
        s164_val_n1 <= s163_val_n1;
    end
    always @(posedge \clk ) begin
        \s165_val  <= \s164_val ;
    end
    always @(posedge \clk ) begin
        s165_val_n1 <= s164_val_n1;
    end
    always @(posedge \clk ) begin
        \s166_val  <= \s165_val ;
    end
    always @(posedge \clk ) begin
        s166_val_n1 <= s165_val_n1;
    end
    always @(posedge \clk ) begin
        \s167_val  <= \s166_val ;
    end
    always @(posedge \clk ) begin
        s167_val_n1 <= s166_val_n1;
    end
    always @(posedge \clk ) begin
        \s168_val  <= \s167_val ;
    end
    always @(posedge \clk ) begin
        s168_val_n1 <= s167_val_n1;
    end
    always @(posedge \clk ) begin
        \s169_val  <= \s168_val ;
    end
    always @(posedge \clk ) begin
        s169_val_n1 <= s168_val_n1;
    end
    always @(posedge \clk ) begin
        \s170_val  <= \s169_val ;
    end
    always @(posedge \clk ) begin
        s170_val_n1 <= s169_val_n1;
    end
    always @(posedge \clk ) begin
        \s171_val  <= \s170_val ;
    end
    always @(posedge \clk ) begin
        s171_val_n1 <= s170_val_n1;
    end
    always @(posedge \clk ) begin
        \s172_val  <= \s171_val ;
    end
    always @(posedge \clk ) begin
        s172_val_n1 <= s171_val_n1;
    end
    always @(posedge \clk ) begin
        \s173_val  <= \s172_val ;
    end
    always @(posedge \clk ) begin
        s173_val_n1 <= s172_val_n1;
    end
    always @(posedge \clk ) begin
        \s174_val  <= \s173_val ;
    end
    always @(posedge \clk ) begin
        s174_val_n1 <= s173_val_n1;
    end
    always @(posedge \clk ) begin
        \s175_val  <= \s174_val ;
    end
    always @(posedge \clk ) begin
        s175_val_n1 <= s174_val_n1;
    end
    always @(posedge \clk ) begin
        \s176_val  <= \s175_val ;
    end
    always @(posedge \clk ) begin
        s176_val_n1 <= s175_val_n1;
    end
    always @(posedge \clk ) begin
        \s177_val  <= \s176_val ;
    end
    always @(posedge \clk ) begin
        s177_val_n1 <= s176_val_n1;
    end
    always @(posedge \clk ) begin
        \s178_val  <= \s177_val ;
    end
    always @(posedge \clk ) begin
        s178_val_n1 <= s177_val_n1;
    end
    always @(posedge \clk ) begin
        \s179_val  <= \s178_val ;
    end
    always @(posedge \clk ) begin
        s179_val_n1 <= s178_val_n1;
    end
    always @(posedge \clk ) begin
        \s180_val  <= \s179_val ;
    end
    always @(posedge \clk ) begin
        s180_val_n1 <= s179_val_n1;
    end
    always @(posedge \clk ) begin
        \s181_val  <= \s180_val ;
    end
    always @(posedge \clk ) begin
        s181_val_n1 <= s180_val_n1;
    end
    always @(posedge \clk ) begin
        \s182_val  <= \s181_val ;
    end
    always @(posedge \clk ) begin
        s182_val_n1 <= s181_val_n1;
    end
    always @(posedge \clk ) begin
        \s183_val  <= \s182_val ;
    end
    always @(posedge \clk ) begin
        s183_val_n1 <= s182_val_n1;
    end
    always @(posedge \clk ) begin
        \s184_val  <= \s183_val ;
    end
    always @(posedge \clk ) begin
        s184_val_n1 <= s183_val_n1;
    end
    always @(posedge \clk ) begin
        \s185_val  <= \s184_val ;
    end
    always @(posedge \clk ) begin
        s185_val_n1 <= s184_val_n1;
    end
    always @(posedge \clk ) begin
        \s186_val  <= \s185_val ;
    end
    always @(posedge \clk ) begin
        s186_val_n1 <= s185_val_n1;
    end
    always @(posedge \clk ) begin
        \s187_val  <= \s186_val ;
    end
    always @(posedge \clk ) begin
        s187_val_n1 <= s186_val_n1;
    end
    always @(posedge \clk ) begin
        \s188_val  <= \s187_val ;
    end
    always @(posedge \clk ) begin
        s188_val_n1 <= s187_val_n1;
    end
    always @(posedge \clk ) begin
        \s189_val  <= \s188_val ;
    end
    always @(posedge \clk ) begin
        s189_val_n1 <= s188_val_n1;
    end
    always @(posedge \clk ) begin
        \s190_val  <= \s189_val ;
    end
    always @(posedge \clk ) begin
        s190_val_n1 <= s189_val_n1;
    end
    always @(posedge \clk ) begin
        \s191_val  <= \s190_val ;
    end
    always @(posedge \clk ) begin
        s191_val_n1 <= s190_val_n1;
    end
    always @(posedge \clk ) begin
        \s192_val  <= \s191_val ;
    end
    always @(posedge \clk ) begin
        s192_val_n1 <= s191_val_n1;
    end
    always @(posedge \clk ) begin
        \s193_val  <= \s192_val ;
    end
    always @(posedge \clk ) begin
        s193_val_n1 <= s192_val_n1;
    end
    always @(posedge \clk ) begin
        \s194_val  <= \s193_val ;
    end
    always @(posedge \clk ) begin
        s194_val_n1 <= s193_val_n1;
    end
    always @(posedge \clk ) begin
        \s195_val  <= \s194_val ;
    end
    always @(posedge \clk ) begin
        s195_val_n1 <= s194_val_n1;
    end
    always @(posedge \clk ) begin
        \s196_val  <= \s195_val ;
    end
    always @(posedge \clk ) begin
        s196_val_n1 <= s195_val_n1;
    end
    always @(posedge \clk ) begin
        \s197_val  <= \s196_val ;
    end
    always @(posedge \clk ) begin
        s197_val_n1 <= s196_val_n1;
    end
    always @(posedge \clk ) begin
        \s198_val  <= \s197_val ;
    end
    always @(posedge \clk ) begin
        s198_val_n1 <= s197_val_n1;
    end
    always @(posedge \clk ) begin
        \s199_val  <= \s198_val ;
    end
    always @(posedge \clk ) begin
        s199_val_n1 <= s198_val_n1;
    end
    always @(posedge \clk ) begin
        \s200_val  <= \s199_val ;
    end
    always @(posedge \clk ) begin
        s200_val_n1 <= s199_val_n1;
    end
    always @(posedge \clk ) begin
        \s201_val  <= \s200_val ;
    end
    always @(posedge \clk ) begin
        s201_val_n1 <= s200_val_n1;
    end
    always @(posedge \clk ) begin
        s201_val_n2 <= val_n2;
    end
    always @(posedge \clk ) begin
        \s202_val  <= \s201_val ;
    end
    always @(posedge \clk ) begin
        s202_val_n1 <= s201_val_n1;
    end
    always @(posedge \clk ) begin
        s202_val_n2 <= s201_val_n2;
    end
    always @(posedge \clk ) begin
        \s203_val  <= \s202_val ;
    end
    always @(posedge \clk ) begin
        s203_val_n1 <= s202_val_n1;
    end
    always @(posedge \clk ) begin
        s203_val_n2 <= s202_val_n2;
    end
    always @(posedge \clk ) begin
        \s204_val  <= \s203_val ;
    end
    always @(posedge \clk ) begin
        s204_val_n1 <= s203_val_n1;
    end
    always @(posedge \clk ) begin
        s204_val_n2 <= s203_val_n2;
    end
    always @(posedge \clk ) begin
        \s205_val  <= \s204_val ;
    end
    always @(posedge \clk ) begin
        s205_val_n1 <= s204_val_n1;
    end
    always @(posedge \clk ) begin
        s205_val_n2 <= s204_val_n2;
    end
    always @(posedge \clk ) begin
        \s206_val  <= \s205_val ;
    end
    always @(posedge \clk ) begin
        s206_val_n1 <= s205_val_n1;
    end
    always @(posedge \clk ) begin
        s206_val_n2 <= s205_val_n2;
    end
    always @(posedge \clk ) begin
        \s207_val  <= \s206_val ;
    end
    always @(posedge \clk ) begin
        s207_val_n1 <= s206_val_n1;
    end
    always @(posedge \clk ) begin
        s207_val_n2 <= s206_val_n2;
    end
    always @(posedge \clk ) begin
        \s208_val  <= \s207_val ;
    end
    always @(posedge \clk ) begin
        s208_val_n1 <= s207_val_n1;
    end
    always @(posedge \clk ) begin
        s208_val_n2 <= s207_val_n2;
    end
    always @(posedge \clk ) begin
        \s209_val  <= \s208_val ;
    end
    always @(posedge \clk ) begin
        s209_val_n1 <= s208_val_n1;
    end
    always @(posedge \clk ) begin
        s209_val_n2 <= s208_val_n2;
    end
    always @(posedge \clk ) begin
        \s210_val  <= \s209_val ;
    end
    always @(posedge \clk ) begin
        s210_val_n1 <= s209_val_n1;
    end
    always @(posedge \clk ) begin
        s210_val_n2 <= s209_val_n2;
    end
    always @(posedge \clk ) begin
        \s211_val  <= \s210_val ;
    end
    always @(posedge \clk ) begin
        s211_val_n1 <= s210_val_n1;
    end
    always @(posedge \clk ) begin
        s211_val_n2 <= s210_val_n2;
    end
    always @(posedge \clk ) begin
        \s212_val  <= \s211_val ;
    end
    always @(posedge \clk ) begin
        s212_val_n1 <= s211_val_n1;
    end
    always @(posedge \clk ) begin
        s212_val_n2 <= s211_val_n2;
    end
    always @(posedge \clk ) begin
        \s213_val  <= \s212_val ;
    end
    always @(posedge \clk ) begin
        s213_val_n1 <= s212_val_n1;
    end
    always @(posedge \clk ) begin
        s213_val_n2 <= s212_val_n2;
    end
    always @(posedge \clk ) begin
        \s214_val  <= \s213_val ;
    end
    always @(posedge \clk ) begin
        s214_val_n1 <= s213_val_n1;
    end
    always @(posedge \clk ) begin
        s214_val_n2 <= s213_val_n2;
    end
    always @(posedge \clk ) begin
        \s215_val  <= \s214_val ;
    end
    always @(posedge \clk ) begin
        s215_val_n1 <= s214_val_n1;
    end
    always @(posedge \clk ) begin
        s215_val_n2 <= s214_val_n2;
    end
    always @(posedge \clk ) begin
        \s216_val  <= \s215_val ;
    end
    always @(posedge \clk ) begin
        s216_val_n1 <= s215_val_n1;
    end
    always @(posedge \clk ) begin
        s216_val_n2 <= s215_val_n2;
    end
    always @(posedge \clk ) begin
        \s217_val  <= \s216_val ;
    end
    always @(posedge \clk ) begin
        s217_val_n1 <= s216_val_n1;
    end
    always @(posedge \clk ) begin
        s217_val_n2 <= s216_val_n2;
    end
    always @(posedge \clk ) begin
        \s218_val  <= \s217_val ;
    end
    always @(posedge \clk ) begin
        s218_val_n1 <= s217_val_n1;
    end
    always @(posedge \clk ) begin
        s218_val_n2 <= s217_val_n2;
    end
    always @(posedge \clk ) begin
        \s219_val  <= \s218_val ;
    end
    always @(posedge \clk ) begin
        s219_val_n1 <= s218_val_n1;
    end
    always @(posedge \clk ) begin
        s219_val_n2 <= s218_val_n2;
    end
    always @(posedge \clk ) begin
        \s220_val  <= \s219_val ;
    end
    always @(posedge \clk ) begin
        s220_val_n1 <= s219_val_n1;
    end
    always @(posedge \clk ) begin
        s220_val_n2 <= s219_val_n2;
    end
    always @(posedge \clk ) begin
        \s221_val  <= \s220_val ;
    end
    always @(posedge \clk ) begin
        s221_val_n1 <= s220_val_n1;
    end
    always @(posedge \clk ) begin
        s221_val_n2 <= s220_val_n2;
    end
    always @(posedge \clk ) begin
        \s222_val  <= \s221_val ;
    end
    always @(posedge \clk ) begin
        s222_val_n1 <= s221_val_n1;
    end
    always @(posedge \clk ) begin
        s222_val_n2 <= s221_val_n2;
    end
    always @(posedge \clk ) begin
        \s223_val  <= \s222_val ;
    end
    always @(posedge \clk ) begin
        s223_val_n1 <= s222_val_n1;
    end
    always @(posedge \clk ) begin
        s223_val_n2 <= s222_val_n2;
    end
    always @(posedge \clk ) begin
        \s224_val  <= \s223_val ;
    end
    always @(posedge \clk ) begin
        s224_val_n1 <= s223_val_n1;
    end
    always @(posedge \clk ) begin
        s224_val_n2 <= s223_val_n2;
    end
    always @(posedge \clk ) begin
        \s225_val  <= \s224_val ;
    end
    always @(posedge \clk ) begin
        s225_val_n1 <= s224_val_n1;
    end
    always @(posedge \clk ) begin
        s225_val_n2 <= s224_val_n2;
    end
    always @(posedge \clk ) begin
        \s226_val  <= \s225_val ;
    end
    always @(posedge \clk ) begin
        s226_val_n1 <= s225_val_n1;
    end
    always @(posedge \clk ) begin
        s226_val_n2 <= s225_val_n2;
    end
    always @(posedge \clk ) begin
        \s227_val  <= \s226_val ;
    end
    always @(posedge \clk ) begin
        s227_val_n1 <= s226_val_n1;
    end
    always @(posedge \clk ) begin
        s227_val_n2 <= s226_val_n2;
    end
    always @(posedge \clk ) begin
        \s228_val  <= \s227_val ;
    end
    always @(posedge \clk ) begin
        s228_val_n1 <= s227_val_n1;
    end
    always @(posedge \clk ) begin
        s228_val_n2 <= s227_val_n2;
    end
    always @(posedge \clk ) begin
        \s229_val  <= \s228_val ;
    end
    always @(posedge \clk ) begin
        s229_val_n1 <= s228_val_n1;
    end
    always @(posedge \clk ) begin
        s229_val_n2 <= s228_val_n2;
    end
    always @(posedge \clk ) begin
        \s230_val  <= \s229_val ;
    end
    always @(posedge \clk ) begin
        s230_val_n1 <= s229_val_n1;
    end
    always @(posedge \clk ) begin
        s230_val_n2 <= s229_val_n2;
    end
    always @(posedge \clk ) begin
        \s231_val  <= \s230_val ;
    end
    always @(posedge \clk ) begin
        s231_val_n1 <= s230_val_n1;
    end
    always @(posedge \clk ) begin
        s231_val_n2 <= s230_val_n2;
    end
    always @(posedge \clk ) begin
        \s232_val  <= \s231_val ;
    end
    always @(posedge \clk ) begin
        s232_val_n1 <= s231_val_n1;
    end
    always @(posedge \clk ) begin
        s232_val_n2 <= s231_val_n2;
    end
    always @(posedge \clk ) begin
        \s233_val  <= \s232_val ;
    end
    always @(posedge \clk ) begin
        s233_val_n1 <= s232_val_n1;
    end
    always @(posedge \clk ) begin
        s233_val_n2 <= s232_val_n2;
    end
    always @(posedge \clk ) begin
        \s234_val  <= \s233_val ;
    end
    always @(posedge \clk ) begin
        s234_val_n1 <= s233_val_n1;
    end
    always @(posedge \clk ) begin
        s234_val_n2 <= s233_val_n2;
    end
    always @(posedge \clk ) begin
        \s235_val  <= \s234_val ;
    end
    always @(posedge \clk ) begin
        s235_val_n1 <= s234_val_n1;
    end
    always @(posedge \clk ) begin
        s235_val_n2 <= s234_val_n2;
    end
    always @(posedge \clk ) begin
        \s236_val  <= \s235_val ;
    end
    always @(posedge \clk ) begin
        s236_val_n1 <= s235_val_n1;
    end
    always @(posedge \clk ) begin
        s236_val_n2 <= s235_val_n2;
    end
    always @(posedge \clk ) begin
        \s237_val  <= \s236_val ;
    end
    always @(posedge \clk ) begin
        s237_val_n1 <= s236_val_n1;
    end
    always @(posedge \clk ) begin
        s237_val_n2 <= s236_val_n2;
    end
    always @(posedge \clk ) begin
        \s238_val  <= \s237_val ;
    end
    always @(posedge \clk ) begin
        s238_val_n1 <= s237_val_n1;
    end
    always @(posedge \clk ) begin
        s238_val_n2 <= s237_val_n2;
    end
    always @(posedge \clk ) begin
        \s239_val  <= \s238_val ;
    end
    always @(posedge \clk ) begin
        s239_val_n1 <= s238_val_n1;
    end
    always @(posedge \clk ) begin
        s239_val_n2 <= s238_val_n2;
    end
    always @(posedge \clk ) begin
        \s240_val  <= \s239_val ;
    end
    always @(posedge \clk ) begin
        s240_val_n1 <= s239_val_n1;
    end
    always @(posedge \clk ) begin
        s240_val_n2 <= s239_val_n2;
    end
    always @(posedge \clk ) begin
        \s241_val  <= \s240_val ;
    end
    always @(posedge \clk ) begin
        s241_val_n1 <= s240_val_n1;
    end
    always @(posedge \clk ) begin
        s241_val_n2 <= s240_val_n2;
    end
    always @(posedge \clk ) begin
        \s242_val  <= \s241_val ;
    end
    always @(posedge \clk ) begin
        s242_val_n1 <= s241_val_n1;
    end
    always @(posedge \clk ) begin
        s242_val_n2 <= s241_val_n2;
    end
    always @(posedge \clk ) begin
        \s243_val  <= \s242_val ;
    end
    always @(posedge \clk ) begin
        s243_val_n1 <= s242_val_n1;
    end
    always @(posedge \clk ) begin
        s243_val_n2 <= s242_val_n2;
    end
    always @(posedge \clk ) begin
        \s244_val  <= \s243_val ;
    end
    always @(posedge \clk ) begin
        s244_val_n1 <= s243_val_n1;
    end
    always @(posedge \clk ) begin
        s244_val_n2 <= s243_val_n2;
    end
    always @(posedge \clk ) begin
        \s245_val  <= \s244_val ;
    end
    always @(posedge \clk ) begin
        s245_val_n1 <= s244_val_n1;
    end
    always @(posedge \clk ) begin
        s245_val_n2 <= s244_val_n2;
    end
    always @(posedge \clk ) begin
        \s246_val  <= \s245_val ;
    end
    always @(posedge \clk ) begin
        s246_val_n1 <= s245_val_n1;
    end
    always @(posedge \clk ) begin
        s246_val_n2 <= s245_val_n2;
    end
    always @(posedge \clk ) begin
        \s247_val  <= \s246_val ;
    end
    always @(posedge \clk ) begin
        s247_val_n1 <= s246_val_n1;
    end
    always @(posedge \clk ) begin
        s247_val_n2 <= s246_val_n2;
    end
    always @(posedge \clk ) begin
        \s248_val  <= \s247_val ;
    end
    always @(posedge \clk ) begin
        s248_val_n1 <= s247_val_n1;
    end
    always @(posedge \clk ) begin
        s248_val_n2 <= s247_val_n2;
    end
    always @(posedge \clk ) begin
        \s249_val  <= \s248_val ;
    end
    always @(posedge \clk ) begin
        s249_val_n1 <= s248_val_n1;
    end
    always @(posedge \clk ) begin
        s249_val_n2 <= s248_val_n2;
    end
    always @(posedge \clk ) begin
        \s250_val  <= \s249_val ;
    end
    always @(posedge \clk ) begin
        s250_val_n1 <= s249_val_n1;
    end
    always @(posedge \clk ) begin
        s250_val_n2 <= s249_val_n2;
    end
    always @(posedge \clk ) begin
        \s251_val  <= \s250_val ;
    end
    always @(posedge \clk ) begin
        s251_val_n1 <= s250_val_n1;
    end
    always @(posedge \clk ) begin
        s251_val_n2 <= s250_val_n2;
    end
    always @(posedge \clk ) begin
        \s252_val  <= \s251_val ;
    end
    always @(posedge \clk ) begin
        s252_val_n1 <= s251_val_n1;
    end
    always @(posedge \clk ) begin
        s252_val_n2 <= s251_val_n2;
    end
    always @(posedge \clk ) begin
        \s253_val  <= \s252_val ;
    end
    always @(posedge \clk ) begin
        s253_val_n1 <= s252_val_n1;
    end
    always @(posedge \clk ) begin
        s253_val_n2 <= s252_val_n2;
    end
    always @(posedge \clk ) begin
        \s254_val  <= \s253_val ;
    end
    always @(posedge \clk ) begin
        s254_val_n1 <= s253_val_n1;
    end
    always @(posedge \clk ) begin
        s254_val_n2 <= s253_val_n2;
    end
    always @(posedge \clk ) begin
        \s255_val  <= \s254_val ;
    end
    always @(posedge \clk ) begin
        s255_val_n1 <= s254_val_n1;
    end
    always @(posedge \clk ) begin
        s255_val_n2 <= s254_val_n2;
    end
    always @(posedge \clk ) begin
        \s256_val  <= \s255_val ;
    end
    always @(posedge \clk ) begin
        s256_val_n1 <= s255_val_n1;
    end
    always @(posedge \clk ) begin
        s256_val_n2 <= s255_val_n2;
    end
    always @(posedge \clk ) begin
        \s257_val  <= \s256_val ;
    end
    always @(posedge \clk ) begin
        s257_val_n1 <= s256_val_n1;
    end
    always @(posedge \clk ) begin
        s257_val_n2 <= s256_val_n2;
    end
    always @(posedge \clk ) begin
        \s258_val  <= \s257_val ;
    end
    always @(posedge \clk ) begin
        s258_val_n1 <= s257_val_n1;
    end
    always @(posedge \clk ) begin
        s258_val_n2 <= s257_val_n2;
    end
    always @(posedge \clk ) begin
        \s259_val  <= \s258_val ;
    end
    always @(posedge \clk ) begin
        s259_val_n1 <= s258_val_n1;
    end
    always @(posedge \clk ) begin
        s259_val_n2 <= s258_val_n2;
    end
    always @(posedge \clk ) begin
        \s260_val  <= \s259_val ;
    end
    always @(posedge \clk ) begin
        s260_val_n1 <= s259_val_n1;
    end
    always @(posedge \clk ) begin
        s260_val_n2 <= s259_val_n2;
    end
    always @(posedge \clk ) begin
        \s261_val  <= \s260_val ;
    end
    always @(posedge \clk ) begin
        s261_val_n1 <= s260_val_n1;
    end
    always @(posedge \clk ) begin
        s261_val_n2 <= s260_val_n2;
    end
    always @(posedge \clk ) begin
        \s262_val  <= \s261_val ;
    end
    always @(posedge \clk ) begin
        s262_val_n1 <= s261_val_n1;
    end
    always @(posedge \clk ) begin
        s262_val_n2 <= s261_val_n2;
    end
    always @(posedge \clk ) begin
        \s263_val  <= \s262_val ;
    end
    always @(posedge \clk ) begin
        s263_val_n1 <= s262_val_n1;
    end
    always @(posedge \clk ) begin
        s263_val_n2 <= s262_val_n2;
    end
    always @(posedge \clk ) begin
        \s264_val  <= \s263_val ;
    end
    always @(posedge \clk ) begin
        s264_val_n1 <= s263_val_n1;
    end
    always @(posedge \clk ) begin
        s264_val_n2 <= s263_val_n2;
    end
    always @(posedge \clk ) begin
        \s265_val  <= \s264_val ;
    end
    always @(posedge \clk ) begin
        s265_val_n1 <= s264_val_n1;
    end
    always @(posedge \clk ) begin
        s265_val_n2 <= s264_val_n2;
    end
    always @(posedge \clk ) begin
        \s266_val  <= \s265_val ;
    end
    always @(posedge \clk ) begin
        s266_val_n1 <= s265_val_n1;
    end
    always @(posedge \clk ) begin
        s266_val_n2 <= s265_val_n2;
    end
    always @(posedge \clk ) begin
        \s267_val  <= \s266_val ;
    end
    always @(posedge \clk ) begin
        s267_val_n1 <= s266_val_n1;
    end
    always @(posedge \clk ) begin
        s267_val_n2 <= s266_val_n2;
    end
    always @(posedge \clk ) begin
        \s268_val  <= \s267_val ;
    end
    always @(posedge \clk ) begin
        s268_val_n1 <= s267_val_n1;
    end
    always @(posedge \clk ) begin
        s268_val_n2 <= s267_val_n2;
    end
    always @(posedge \clk ) begin
        \s269_val  <= \s268_val ;
    end
    always @(posedge \clk ) begin
        s269_val_n1 <= s268_val_n1;
    end
    always @(posedge \clk ) begin
        s269_val_n2 <= s268_val_n2;
    end
    always @(posedge \clk ) begin
        \s270_val  <= \s269_val ;
    end
    always @(posedge \clk ) begin
        s270_val_n1 <= s269_val_n1;
    end
    always @(posedge \clk ) begin
        s270_val_n2 <= s269_val_n2;
    end
    always @(posedge \clk ) begin
        \s271_val  <= \s270_val ;
    end
    always @(posedge \clk ) begin
        s271_val_n1 <= s270_val_n1;
    end
    always @(posedge \clk ) begin
        s271_val_n2 <= s270_val_n2;
    end
    always @(posedge \clk ) begin
        \s272_val  <= \s271_val ;
    end
    always @(posedge \clk ) begin
        s272_val_n1 <= s271_val_n1;
    end
    always @(posedge \clk ) begin
        s272_val_n2 <= s271_val_n2;
    end
    always @(posedge \clk ) begin
        \s273_val  <= \s272_val ;
    end
    always @(posedge \clk ) begin
        s273_val_n1 <= s272_val_n1;
    end
    always @(posedge \clk ) begin
        s273_val_n2 <= s272_val_n2;
    end
    always @(posedge \clk ) begin
        \s274_val  <= \s273_val ;
    end
    always @(posedge \clk ) begin
        s274_val_n1 <= s273_val_n1;
    end
    always @(posedge \clk ) begin
        s274_val_n2 <= s273_val_n2;
    end
    always @(posedge \clk ) begin
        \s275_val  <= \s274_val ;
    end
    always @(posedge \clk ) begin
        s275_val_n1 <= s274_val_n1;
    end
    always @(posedge \clk ) begin
        s275_val_n2 <= s274_val_n2;
    end
    always @(posedge \clk ) begin
        \s276_val  <= \s275_val ;
    end
    always @(posedge \clk ) begin
        s276_val_n1 <= s275_val_n1;
    end
    always @(posedge \clk ) begin
        s276_val_n2 <= s275_val_n2;
    end
    always @(posedge \clk ) begin
        \s277_val  <= \s276_val ;
    end
    always @(posedge \clk ) begin
        s277_val_n1 <= s276_val_n1;
    end
    always @(posedge \clk ) begin
        s277_val_n2 <= s276_val_n2;
    end
    always @(posedge \clk ) begin
        \s278_val  <= \s277_val ;
    end
    always @(posedge \clk ) begin
        s278_val_n1 <= s277_val_n1;
    end
    always @(posedge \clk ) begin
        s278_val_n2 <= s277_val_n2;
    end
    always @(posedge \clk ) begin
        \s279_val  <= \s278_val ;
    end
    always @(posedge \clk ) begin
        s279_val_n1 <= s278_val_n1;
    end
    always @(posedge \clk ) begin
        s279_val_n2 <= s278_val_n2;
    end
    always @(posedge \clk ) begin
        \s280_val  <= \s279_val ;
    end
    always @(posedge \clk ) begin
        s280_val_n1 <= s279_val_n1;
    end
    always @(posedge \clk ) begin
        s280_val_n2 <= s279_val_n2;
    end
    always @(posedge \clk ) begin
        \s281_val  <= \s280_val ;
    end
    always @(posedge \clk ) begin
        s281_val_n1 <= s280_val_n1;
    end
    always @(posedge \clk ) begin
        s281_val_n2 <= s280_val_n2;
    end
    always @(posedge \clk ) begin
        \s282_val  <= \s281_val ;
    end
    always @(posedge \clk ) begin
        s282_val_n1 <= s281_val_n1;
    end
    always @(posedge \clk ) begin
        s282_val_n2 <= s281_val_n2;
    end
    always @(posedge \clk ) begin
        \s283_val  <= \s282_val ;
    end
    always @(posedge \clk ) begin
        s283_val_n1 <= s282_val_n1;
    end
    always @(posedge \clk ) begin
        s283_val_n2 <= s282_val_n2;
    end
    always @(posedge \clk ) begin
        \s284_val  <= \s283_val ;
    end
    always @(posedge \clk ) begin
        s284_val_n1 <= s283_val_n1;
    end
    always @(posedge \clk ) begin
        s284_val_n2 <= s283_val_n2;
    end
    always @(posedge \clk ) begin
        \s285_val  <= \s284_val ;
    end
    always @(posedge \clk ) begin
        s285_val_n1 <= s284_val_n1;
    end
    always @(posedge \clk ) begin
        s285_val_n2 <= s284_val_n2;
    end
    always @(posedge \clk ) begin
        \s286_val  <= \s285_val ;
    end
    always @(posedge \clk ) begin
        s286_val_n1 <= s285_val_n1;
    end
    always @(posedge \clk ) begin
        s286_val_n2 <= s285_val_n2;
    end
    always @(posedge \clk ) begin
        \s287_val  <= \s286_val ;
    end
    always @(posedge \clk ) begin
        s287_val_n1 <= s286_val_n1;
    end
    always @(posedge \clk ) begin
        s287_val_n2 <= s286_val_n2;
    end
    always @(posedge \clk ) begin
        \s288_val  <= \s287_val ;
    end
    always @(posedge \clk ) begin
        s288_val_n1 <= s287_val_n1;
    end
    always @(posedge \clk ) begin
        s288_val_n2 <= s287_val_n2;
    end
    always @(posedge \clk ) begin
        \s289_val  <= \s288_val ;
    end
    always @(posedge \clk ) begin
        s289_val_n1 <= s288_val_n1;
    end
    always @(posedge \clk ) begin
        s289_val_n2 <= s288_val_n2;
    end
    always @(posedge \clk ) begin
        \s290_val  <= \s289_val ;
    end
    always @(posedge \clk ) begin
        s290_val_n1 <= s289_val_n1;
    end
    always @(posedge \clk ) begin
        s290_val_n2 <= s289_val_n2;
    end
    always @(posedge \clk ) begin
        \s291_val  <= \s290_val ;
    end
    always @(posedge \clk ) begin
        s291_val_n1 <= s290_val_n1;
    end
    always @(posedge \clk ) begin
        s291_val_n2 <= s290_val_n2;
    end
    always @(posedge \clk ) begin
        \s292_val  <= \s291_val ;
    end
    always @(posedge \clk ) begin
        s292_val_n1 <= s291_val_n1;
    end
    always @(posedge \clk ) begin
        s292_val_n2 <= s291_val_n2;
    end
    always @(posedge \clk ) begin
        \s293_val  <= \s292_val ;
    end
    always @(posedge \clk ) begin
        s293_val_n1 <= s292_val_n1;
    end
    always @(posedge \clk ) begin
        s293_val_n2 <= s292_val_n2;
    end
    always @(posedge \clk ) begin
        \s294_val  <= \s293_val ;
    end
    always @(posedge \clk ) begin
        s294_val_n1 <= s293_val_n1;
    end
    always @(posedge \clk ) begin
        s294_val_n2 <= s293_val_n2;
    end
    always @(posedge \clk ) begin
        \s295_val  <= \s294_val ;
    end
    always @(posedge \clk ) begin
        s295_val_n1 <= s294_val_n1;
    end
    always @(posedge \clk ) begin
        s295_val_n2 <= s294_val_n2;
    end
    always @(posedge \clk ) begin
        \s296_val  <= \s295_val ;
    end
    always @(posedge \clk ) begin
        s296_val_n1 <= s295_val_n1;
    end
    always @(posedge \clk ) begin
        s296_val_n2 <= s295_val_n2;
    end
    always @(posedge \clk ) begin
        \s297_val  <= \s296_val ;
    end
    always @(posedge \clk ) begin
        s297_val_n1 <= s296_val_n1;
    end
    always @(posedge \clk ) begin
        s297_val_n2 <= s296_val_n2;
    end
    always @(posedge \clk ) begin
        \s298_val  <= \s297_val ;
    end
    always @(posedge \clk ) begin
        s298_val_n1 <= s297_val_n1;
    end
    always @(posedge \clk ) begin
        s298_val_n2 <= s297_val_n2;
    end
    always @(posedge \clk ) begin
        \s299_val  <= \s298_val ;
    end
    always @(posedge \clk ) begin
        s299_val_n1 <= s298_val_n1;
    end
    always @(posedge \clk ) begin
        s299_val_n2 <= s298_val_n2;
    end
    always @(posedge \clk ) begin
        \s300_val  <= \s299_val ;
    end
    always @(posedge \clk ) begin
        s300_val_n1 <= s299_val_n1;
    end
    always @(posedge \clk ) begin
        s300_val_n2 <= s299_val_n2;
    end
    always @(posedge \clk ) begin
        \s301_val  <= \s300_val ;
    end
    always @(posedge \clk ) begin
        s301_val_n1 <= s300_val_n1;
    end
    always @(posedge \clk ) begin
        s301_val_n2 <= s300_val_n2;
    end
    always @(posedge \clk ) begin
        s301_val_n3 <= val_n3;
    end
    always @(posedge \clk ) begin
        \s302_val  <= \s301_val ;
    end
    always @(posedge \clk ) begin
        s302_val_n1 <= s301_val_n1;
    end
    always @(posedge \clk ) begin
        s302_val_n2 <= s301_val_n2;
    end
    always @(posedge \clk ) begin
        s302_val_n3 <= s301_val_n3;
    end
    always @(posedge \clk ) begin
        \s303_val  <= \s302_val ;
    end
    always @(posedge \clk ) begin
        s303_val_n1 <= s302_val_n1;
    end
    always @(posedge \clk ) begin
        s303_val_n2 <= s302_val_n2;
    end
    always @(posedge \clk ) begin
        s303_val_n3 <= s302_val_n3;
    end
    always @(posedge \clk ) begin
        \s304_val  <= \s303_val ;
    end
    always @(posedge \clk ) begin
        s304_val_n1 <= s303_val_n1;
    end
    always @(posedge \clk ) begin
        s304_val_n2 <= s303_val_n2;
    end
    always @(posedge \clk ) begin
        s304_val_n3 <= s303_val_n3;
    end
    always @(posedge \clk ) begin
        \s305_val  <= \s304_val ;
    end
    always @(posedge \clk ) begin
        s305_val_n1 <= s304_val_n1;
    end
    always @(posedge \clk ) begin
        s305_val_n2 <= s304_val_n2;
    end
    always @(posedge \clk ) begin
        s305_val_n3 <= s304_val_n3;
    end
    always @(posedge \clk ) begin
        \s306_val  <= \s305_val ;
    end
    always @(posedge \clk ) begin
        s306_val_n1 <= s305_val_n1;
    end
    always @(posedge \clk ) begin
        s306_val_n2 <= s305_val_n2;
    end
    always @(posedge \clk ) begin
        s306_val_n3 <= s305_val_n3;
    end
    always @(posedge \clk ) begin
        \s307_val  <= \s306_val ;
    end
    always @(posedge \clk ) begin
        s307_val_n1 <= s306_val_n1;
    end
    always @(posedge \clk ) begin
        s307_val_n2 <= s306_val_n2;
    end
    always @(posedge \clk ) begin
        s307_val_n3 <= s306_val_n3;
    end
    always @(posedge \clk ) begin
        \s308_val  <= \s307_val ;
    end
    always @(posedge \clk ) begin
        s308_val_n1 <= s307_val_n1;
    end
    always @(posedge \clk ) begin
        s308_val_n2 <= s307_val_n2;
    end
    always @(posedge \clk ) begin
        s308_val_n3 <= s307_val_n3;
    end
    always @(posedge \clk ) begin
        \s309_val  <= \s308_val ;
    end
    always @(posedge \clk ) begin
        s309_val_n1 <= s308_val_n1;
    end
    always @(posedge \clk ) begin
        s309_val_n2 <= s308_val_n2;
    end
    always @(posedge \clk ) begin
        s309_val_n3 <= s308_val_n3;
    end
    always @(posedge \clk ) begin
        \s310_val  <= \s309_val ;
    end
    always @(posedge \clk ) begin
        s310_val_n1 <= s309_val_n1;
    end
    always @(posedge \clk ) begin
        s310_val_n2 <= s309_val_n2;
    end
    always @(posedge \clk ) begin
        s310_val_n3 <= s309_val_n3;
    end
    always @(posedge \clk ) begin
        \s311_val  <= \s310_val ;
    end
    always @(posedge \clk ) begin
        s311_val_n1 <= s310_val_n1;
    end
    always @(posedge \clk ) begin
        s311_val_n2 <= s310_val_n2;
    end
    always @(posedge \clk ) begin
        s311_val_n3 <= s310_val_n3;
    end
    always @(posedge \clk ) begin
        \s312_val  <= \s311_val ;
    end
    always @(posedge \clk ) begin
        s312_val_n1 <= s311_val_n1;
    end
    always @(posedge \clk ) begin
        s312_val_n2 <= s311_val_n2;
    end
    always @(posedge \clk ) begin
        s312_val_n3 <= s311_val_n3;
    end
    always @(posedge \clk ) begin
        \s313_val  <= \s312_val ;
    end
    always @(posedge \clk ) begin
        s313_val_n1 <= s312_val_n1;
    end
    always @(posedge \clk ) begin
        s313_val_n2 <= s312_val_n2;
    end
    always @(posedge \clk ) begin
        s313_val_n3 <= s312_val_n3;
    end
    always @(posedge \clk ) begin
        \s314_val  <= \s313_val ;
    end
    always @(posedge \clk ) begin
        s314_val_n1 <= s313_val_n1;
    end
    always @(posedge \clk ) begin
        s314_val_n2 <= s313_val_n2;
    end
    always @(posedge \clk ) begin
        s314_val_n3 <= s313_val_n3;
    end
    always @(posedge \clk ) begin
        \s315_val  <= \s314_val ;
    end
    always @(posedge \clk ) begin
        s315_val_n1 <= s314_val_n1;
    end
    always @(posedge \clk ) begin
        s315_val_n2 <= s314_val_n2;
    end
    always @(posedge \clk ) begin
        s315_val_n3 <= s314_val_n3;
    end
    always @(posedge \clk ) begin
        \s316_val  <= \s315_val ;
    end
    always @(posedge \clk ) begin
        s316_val_n1 <= s315_val_n1;
    end
    always @(posedge \clk ) begin
        s316_val_n2 <= s315_val_n2;
    end
    always @(posedge \clk ) begin
        s316_val_n3 <= s315_val_n3;
    end
    always @(posedge \clk ) begin
        \s317_val  <= \s316_val ;
    end
    always @(posedge \clk ) begin
        s317_val_n1 <= s316_val_n1;
    end
    always @(posedge \clk ) begin
        s317_val_n2 <= s316_val_n2;
    end
    always @(posedge \clk ) begin
        s317_val_n3 <= s316_val_n3;
    end
    always @(posedge \clk ) begin
        \s318_val  <= \s317_val ;
    end
    always @(posedge \clk ) begin
        s318_val_n1 <= s317_val_n1;
    end
    always @(posedge \clk ) begin
        s318_val_n2 <= s317_val_n2;
    end
    always @(posedge \clk ) begin
        s318_val_n3 <= s317_val_n3;
    end
    always @(posedge \clk ) begin
        \s319_val  <= \s318_val ;
    end
    always @(posedge \clk ) begin
        s319_val_n1 <= s318_val_n1;
    end
    always @(posedge \clk ) begin
        s319_val_n2 <= s318_val_n2;
    end
    always @(posedge \clk ) begin
        s319_val_n3 <= s318_val_n3;
    end
    always @(posedge \clk ) begin
        \s320_val  <= \s319_val ;
    end
    always @(posedge \clk ) begin
        s320_val_n1 <= s319_val_n1;
    end
    always @(posedge \clk ) begin
        s320_val_n2 <= s319_val_n2;
    end
    always @(posedge \clk ) begin
        s320_val_n3 <= s319_val_n3;
    end
    always @(posedge \clk ) begin
        \s321_val  <= \s320_val ;
    end
    always @(posedge \clk ) begin
        s321_val_n1 <= s320_val_n1;
    end
    always @(posedge \clk ) begin
        s321_val_n2 <= s320_val_n2;
    end
    always @(posedge \clk ) begin
        s321_val_n3 <= s320_val_n3;
    end
    always @(posedge \clk ) begin
        \s322_val  <= \s321_val ;
    end
    always @(posedge \clk ) begin
        s322_val_n1 <= s321_val_n1;
    end
    always @(posedge \clk ) begin
        s322_val_n2 <= s321_val_n2;
    end
    always @(posedge \clk ) begin
        s322_val_n3 <= s321_val_n3;
    end
    always @(posedge \clk ) begin
        \s323_val  <= \s322_val ;
    end
    always @(posedge \clk ) begin
        s323_val_n1 <= s322_val_n1;
    end
    always @(posedge \clk ) begin
        s323_val_n2 <= s322_val_n2;
    end
    always @(posedge \clk ) begin
        s323_val_n3 <= s322_val_n3;
    end
    always @(posedge \clk ) begin
        \s324_val  <= \s323_val ;
    end
    always @(posedge \clk ) begin
        s324_val_n1 <= s323_val_n1;
    end
    always @(posedge \clk ) begin
        s324_val_n2 <= s323_val_n2;
    end
    always @(posedge \clk ) begin
        s324_val_n3 <= s323_val_n3;
    end
    always @(posedge \clk ) begin
        \s325_val  <= \s324_val ;
    end
    always @(posedge \clk ) begin
        s325_val_n1 <= s324_val_n1;
    end
    always @(posedge \clk ) begin
        s325_val_n2 <= s324_val_n2;
    end
    always @(posedge \clk ) begin
        s325_val_n3 <= s324_val_n3;
    end
    always @(posedge \clk ) begin
        \s326_val  <= \s325_val ;
    end
    always @(posedge \clk ) begin
        s326_val_n1 <= s325_val_n1;
    end
    always @(posedge \clk ) begin
        s326_val_n2 <= s325_val_n2;
    end
    always @(posedge \clk ) begin
        s326_val_n3 <= s325_val_n3;
    end
    always @(posedge \clk ) begin
        \s327_val  <= \s326_val ;
    end
    always @(posedge \clk ) begin
        s327_val_n1 <= s326_val_n1;
    end
    always @(posedge \clk ) begin
        s327_val_n2 <= s326_val_n2;
    end
    always @(posedge \clk ) begin
        s327_val_n3 <= s326_val_n3;
    end
    always @(posedge \clk ) begin
        \s328_val  <= \s327_val ;
    end
    always @(posedge \clk ) begin
        s328_val_n1 <= s327_val_n1;
    end
    always @(posedge \clk ) begin
        s328_val_n2 <= s327_val_n2;
    end
    always @(posedge \clk ) begin
        s328_val_n3 <= s327_val_n3;
    end
    always @(posedge \clk ) begin
        \s329_val  <= \s328_val ;
    end
    always @(posedge \clk ) begin
        s329_val_n1 <= s328_val_n1;
    end
    always @(posedge \clk ) begin
        s329_val_n2 <= s328_val_n2;
    end
    always @(posedge \clk ) begin
        s329_val_n3 <= s328_val_n3;
    end
    always @(posedge \clk ) begin
        \s330_val  <= \s329_val ;
    end
    always @(posedge \clk ) begin
        s330_val_n1 <= s329_val_n1;
    end
    always @(posedge \clk ) begin
        s330_val_n2 <= s329_val_n2;
    end
    always @(posedge \clk ) begin
        s330_val_n3 <= s329_val_n3;
    end
    always @(posedge \clk ) begin
        \s331_val  <= \s330_val ;
    end
    always @(posedge \clk ) begin
        s331_val_n1 <= s330_val_n1;
    end
    always @(posedge \clk ) begin
        s331_val_n2 <= s330_val_n2;
    end
    always @(posedge \clk ) begin
        s331_val_n3 <= s330_val_n3;
    end
    always @(posedge \clk ) begin
        \s332_val  <= \s331_val ;
    end
    always @(posedge \clk ) begin
        s332_val_n1 <= s331_val_n1;
    end
    always @(posedge \clk ) begin
        s332_val_n2 <= s331_val_n2;
    end
    always @(posedge \clk ) begin
        s332_val_n3 <= s331_val_n3;
    end
    always @(posedge \clk ) begin
        \s333_val  <= \s332_val ;
    end
    always @(posedge \clk ) begin
        s333_val_n1 <= s332_val_n1;
    end
    always @(posedge \clk ) begin
        s333_val_n2 <= s332_val_n2;
    end
    always @(posedge \clk ) begin
        s333_val_n3 <= s332_val_n3;
    end
    always @(posedge \clk ) begin
        \s334_val  <= \s333_val ;
    end
    always @(posedge \clk ) begin
        s334_val_n1 <= s333_val_n1;
    end
    always @(posedge \clk ) begin
        s334_val_n2 <= s333_val_n2;
    end
    always @(posedge \clk ) begin
        s334_val_n3 <= s333_val_n3;
    end
    always @(posedge \clk ) begin
        \s335_val  <= \s334_val ;
    end
    always @(posedge \clk ) begin
        s335_val_n1 <= s334_val_n1;
    end
    always @(posedge \clk ) begin
        s335_val_n2 <= s334_val_n2;
    end
    always @(posedge \clk ) begin
        s335_val_n3 <= s334_val_n3;
    end
    always @(posedge \clk ) begin
        \s336_val  <= \s335_val ;
    end
    always @(posedge \clk ) begin
        s336_val_n1 <= s335_val_n1;
    end
    always @(posedge \clk ) begin
        s336_val_n2 <= s335_val_n2;
    end
    always @(posedge \clk ) begin
        s336_val_n3 <= s335_val_n3;
    end
    always @(posedge \clk ) begin
        \s337_val  <= \s336_val ;
    end
    always @(posedge \clk ) begin
        s337_val_n1 <= s336_val_n1;
    end
    always @(posedge \clk ) begin
        s337_val_n2 <= s336_val_n2;
    end
    always @(posedge \clk ) begin
        s337_val_n3 <= s336_val_n3;
    end
    always @(posedge \clk ) begin
        \s338_val  <= \s337_val ;
    end
    always @(posedge \clk ) begin
        s338_val_n1 <= s337_val_n1;
    end
    always @(posedge \clk ) begin
        s338_val_n2 <= s337_val_n2;
    end
    always @(posedge \clk ) begin
        s338_val_n3 <= s337_val_n3;
    end
    always @(posedge \clk ) begin
        \s339_val  <= \s338_val ;
    end
    always @(posedge \clk ) begin
        s339_val_n1 <= s338_val_n1;
    end
    always @(posedge \clk ) begin
        s339_val_n2 <= s338_val_n2;
    end
    always @(posedge \clk ) begin
        s339_val_n3 <= s338_val_n3;
    end
    always @(posedge \clk ) begin
        \s340_val  <= \s339_val ;
    end
    always @(posedge \clk ) begin
        s340_val_n1 <= s339_val_n1;
    end
    always @(posedge \clk ) begin
        s340_val_n2 <= s339_val_n2;
    end
    always @(posedge \clk ) begin
        s340_val_n3 <= s339_val_n3;
    end
    always @(posedge \clk ) begin
        \s341_val  <= \s340_val ;
    end
    always @(posedge \clk ) begin
        s341_val_n1 <= s340_val_n1;
    end
    always @(posedge \clk ) begin
        s341_val_n2 <= s340_val_n2;
    end
    always @(posedge \clk ) begin
        s341_val_n3 <= s340_val_n3;
    end
    always @(posedge \clk ) begin
        \s342_val  <= \s341_val ;
    end
    always @(posedge \clk ) begin
        s342_val_n1 <= s341_val_n1;
    end
    always @(posedge \clk ) begin
        s342_val_n2 <= s341_val_n2;
    end
    always @(posedge \clk ) begin
        s342_val_n3 <= s341_val_n3;
    end
    always @(posedge \clk ) begin
        \s343_val  <= \s342_val ;
    end
    always @(posedge \clk ) begin
        s343_val_n1 <= s342_val_n1;
    end
    always @(posedge \clk ) begin
        s343_val_n2 <= s342_val_n2;
    end
    always @(posedge \clk ) begin
        s343_val_n3 <= s342_val_n3;
    end
    always @(posedge \clk ) begin
        \s344_val  <= \s343_val ;
    end
    always @(posedge \clk ) begin
        s344_val_n1 <= s343_val_n1;
    end
    always @(posedge \clk ) begin
        s344_val_n2 <= s343_val_n2;
    end
    always @(posedge \clk ) begin
        s344_val_n3 <= s343_val_n3;
    end
    always @(posedge \clk ) begin
        \s345_val  <= \s344_val ;
    end
    always @(posedge \clk ) begin
        s345_val_n1 <= s344_val_n1;
    end
    always @(posedge \clk ) begin
        s345_val_n2 <= s344_val_n2;
    end
    always @(posedge \clk ) begin
        s345_val_n3 <= s344_val_n3;
    end
    always @(posedge \clk ) begin
        \s346_val  <= \s345_val ;
    end
    always @(posedge \clk ) begin
        s346_val_n1 <= s345_val_n1;
    end
    always @(posedge \clk ) begin
        s346_val_n2 <= s345_val_n2;
    end
    always @(posedge \clk ) begin
        s346_val_n3 <= s345_val_n3;
    end
    always @(posedge \clk ) begin
        \s347_val  <= \s346_val ;
    end
    always @(posedge \clk ) begin
        s347_val_n1 <= s346_val_n1;
    end
    always @(posedge \clk ) begin
        s347_val_n2 <= s346_val_n2;
    end
    always @(posedge \clk ) begin
        s347_val_n3 <= s346_val_n3;
    end
    always @(posedge \clk ) begin
        \s348_val  <= \s347_val ;
    end
    always @(posedge \clk ) begin
        s348_val_n1 <= s347_val_n1;
    end
    always @(posedge \clk ) begin
        s348_val_n2 <= s347_val_n2;
    end
    always @(posedge \clk ) begin
        s348_val_n3 <= s347_val_n3;
    end
    always @(posedge \clk ) begin
        \s349_val  <= \s348_val ;
    end
    always @(posedge \clk ) begin
        s349_val_n1 <= s348_val_n1;
    end
    always @(posedge \clk ) begin
        s349_val_n2 <= s348_val_n2;
    end
    always @(posedge \clk ) begin
        s349_val_n3 <= s348_val_n3;
    end
    always @(posedge \clk ) begin
        \s350_val  <= \s349_val ;
    end
    always @(posedge \clk ) begin
        s350_val_n1 <= s349_val_n1;
    end
    always @(posedge \clk ) begin
        s350_val_n2 <= s349_val_n2;
    end
    always @(posedge \clk ) begin
        s350_val_n3 <= s349_val_n3;
    end
    always @(posedge \clk ) begin
        \s351_val  <= \s350_val ;
    end
    always @(posedge \clk ) begin
        s351_val_n1 <= s350_val_n1;
    end
    always @(posedge \clk ) begin
        s351_val_n2 <= s350_val_n2;
    end
    always @(posedge \clk ) begin
        s351_val_n3 <= s350_val_n3;
    end
    always @(posedge \clk ) begin
        \s352_val  <= \s351_val ;
    end
    always @(posedge \clk ) begin
        s352_val_n1 <= s351_val_n1;
    end
    always @(posedge \clk ) begin
        s352_val_n2 <= s351_val_n2;
    end
    always @(posedge \clk ) begin
        s352_val_n3 <= s351_val_n3;
    end
    always @(posedge \clk ) begin
        \s353_val  <= \s352_val ;
    end
    always @(posedge \clk ) begin
        s353_val_n1 <= s352_val_n1;
    end
    always @(posedge \clk ) begin
        s353_val_n2 <= s352_val_n2;
    end
    always @(posedge \clk ) begin
        s353_val_n3 <= s352_val_n3;
    end
    always @(posedge \clk ) begin
        \s354_val  <= \s353_val ;
    end
    always @(posedge \clk ) begin
        s354_val_n1 <= s353_val_n1;
    end
    always @(posedge \clk ) begin
        s354_val_n2 <= s353_val_n2;
    end
    always @(posedge \clk ) begin
        s354_val_n3 <= s353_val_n3;
    end
    always @(posedge \clk ) begin
        \s355_val  <= \s354_val ;
    end
    always @(posedge \clk ) begin
        s355_val_n1 <= s354_val_n1;
    end
    always @(posedge \clk ) begin
        s355_val_n2 <= s354_val_n2;
    end
    always @(posedge \clk ) begin
        s355_val_n3 <= s354_val_n3;
    end
    always @(posedge \clk ) begin
        \s356_val  <= \s355_val ;
    end
    always @(posedge \clk ) begin
        s356_val_n1 <= s355_val_n1;
    end
    always @(posedge \clk ) begin
        s356_val_n2 <= s355_val_n2;
    end
    always @(posedge \clk ) begin
        s356_val_n3 <= s355_val_n3;
    end
    always @(posedge \clk ) begin
        \s357_val  <= \s356_val ;
    end
    always @(posedge \clk ) begin
        s357_val_n1 <= s356_val_n1;
    end
    always @(posedge \clk ) begin
        s357_val_n2 <= s356_val_n2;
    end
    always @(posedge \clk ) begin
        s357_val_n3 <= s356_val_n3;
    end
    always @(posedge \clk ) begin
        \s358_val  <= \s357_val ;
    end
    always @(posedge \clk ) begin
        s358_val_n1 <= s357_val_n1;
    end
    always @(posedge \clk ) begin
        s358_val_n2 <= s357_val_n2;
    end
    always @(posedge \clk ) begin
        s358_val_n3 <= s357_val_n3;
    end
    always @(posedge \clk ) begin
        \s359_val  <= \s358_val ;
    end
    always @(posedge \clk ) begin
        s359_val_n1 <= s358_val_n1;
    end
    always @(posedge \clk ) begin
        s359_val_n2 <= s358_val_n2;
    end
    always @(posedge \clk ) begin
        s359_val_n3 <= s358_val_n3;
    end
    always @(posedge \clk ) begin
        \s360_val  <= \s359_val ;
    end
    always @(posedge \clk ) begin
        s360_val_n1 <= s359_val_n1;
    end
    always @(posedge \clk ) begin
        s360_val_n2 <= s359_val_n2;
    end
    always @(posedge \clk ) begin
        s360_val_n3 <= s359_val_n3;
    end
    always @(posedge \clk ) begin
        \s361_val  <= \s360_val ;
    end
    always @(posedge \clk ) begin
        s361_val_n1 <= s360_val_n1;
    end
    always @(posedge \clk ) begin
        s361_val_n2 <= s360_val_n2;
    end
    always @(posedge \clk ) begin
        s361_val_n3 <= s360_val_n3;
    end
    always @(posedge \clk ) begin
        \s362_val  <= \s361_val ;
    end
    always @(posedge \clk ) begin
        s362_val_n1 <= s361_val_n1;
    end
    always @(posedge \clk ) begin
        s362_val_n2 <= s361_val_n2;
    end
    always @(posedge \clk ) begin
        s362_val_n3 <= s361_val_n3;
    end
    always @(posedge \clk ) begin
        \s363_val  <= \s362_val ;
    end
    always @(posedge \clk ) begin
        s363_val_n1 <= s362_val_n1;
    end
    always @(posedge \clk ) begin
        s363_val_n2 <= s362_val_n2;
    end
    always @(posedge \clk ) begin
        s363_val_n3 <= s362_val_n3;
    end
    always @(posedge \clk ) begin
        \s364_val  <= \s363_val ;
    end
    always @(posedge \clk ) begin
        s364_val_n1 <= s363_val_n1;
    end
    always @(posedge \clk ) begin
        s364_val_n2 <= s363_val_n2;
    end
    always @(posedge \clk ) begin
        s364_val_n3 <= s363_val_n3;
    end
    always @(posedge \clk ) begin
        \s365_val  <= \s364_val ;
    end
    always @(posedge \clk ) begin
        s365_val_n1 <= s364_val_n1;
    end
    always @(posedge \clk ) begin
        s365_val_n2 <= s364_val_n2;
    end
    always @(posedge \clk ) begin
        s365_val_n3 <= s364_val_n3;
    end
    always @(posedge \clk ) begin
        \s366_val  <= \s365_val ;
    end
    always @(posedge \clk ) begin
        s366_val_n1 <= s365_val_n1;
    end
    always @(posedge \clk ) begin
        s366_val_n2 <= s365_val_n2;
    end
    always @(posedge \clk ) begin
        s366_val_n3 <= s365_val_n3;
    end
    always @(posedge \clk ) begin
        \s367_val  <= \s366_val ;
    end
    always @(posedge \clk ) begin
        s367_val_n1 <= s366_val_n1;
    end
    always @(posedge \clk ) begin
        s367_val_n2 <= s366_val_n2;
    end
    always @(posedge \clk ) begin
        s367_val_n3 <= s366_val_n3;
    end
    always @(posedge \clk ) begin
        \s368_val  <= \s367_val ;
    end
    always @(posedge \clk ) begin
        s368_val_n1 <= s367_val_n1;
    end
    always @(posedge \clk ) begin
        s368_val_n2 <= s367_val_n2;
    end
    always @(posedge \clk ) begin
        s368_val_n3 <= s367_val_n3;
    end
    always @(posedge \clk ) begin
        \s369_val  <= \s368_val ;
    end
    always @(posedge \clk ) begin
        s369_val_n1 <= s368_val_n1;
    end
    always @(posedge \clk ) begin
        s369_val_n2 <= s368_val_n2;
    end
    always @(posedge \clk ) begin
        s369_val_n3 <= s368_val_n3;
    end
    always @(posedge \clk ) begin
        \s370_val  <= \s369_val ;
    end
    always @(posedge \clk ) begin
        s370_val_n1 <= s369_val_n1;
    end
    always @(posedge \clk ) begin
        s370_val_n2 <= s369_val_n2;
    end
    always @(posedge \clk ) begin
        s370_val_n3 <= s369_val_n3;
    end
    always @(posedge \clk ) begin
        \s371_val  <= \s370_val ;
    end
    always @(posedge \clk ) begin
        s371_val_n1 <= s370_val_n1;
    end
    always @(posedge \clk ) begin
        s371_val_n2 <= s370_val_n2;
    end
    always @(posedge \clk ) begin
        s371_val_n3 <= s370_val_n3;
    end
    always @(posedge \clk ) begin
        \s372_val  <= \s371_val ;
    end
    always @(posedge \clk ) begin
        s372_val_n1 <= s371_val_n1;
    end
    always @(posedge \clk ) begin
        s372_val_n2 <= s371_val_n2;
    end
    always @(posedge \clk ) begin
        s372_val_n3 <= s371_val_n3;
    end
    always @(posedge \clk ) begin
        \s373_val  <= \s372_val ;
    end
    always @(posedge \clk ) begin
        s373_val_n1 <= s372_val_n1;
    end
    always @(posedge \clk ) begin
        s373_val_n2 <= s372_val_n2;
    end
    always @(posedge \clk ) begin
        s373_val_n3 <= s372_val_n3;
    end
    always @(posedge \clk ) begin
        \s374_val  <= \s373_val ;
    end
    always @(posedge \clk ) begin
        s374_val_n1 <= s373_val_n1;
    end
    always @(posedge \clk ) begin
        s374_val_n2 <= s373_val_n2;
    end
    always @(posedge \clk ) begin
        s374_val_n3 <= s373_val_n3;
    end
    always @(posedge \clk ) begin
        \s375_val  <= \s374_val ;
    end
    always @(posedge \clk ) begin
        s375_val_n1 <= s374_val_n1;
    end
    always @(posedge \clk ) begin
        s375_val_n2 <= s374_val_n2;
    end
    always @(posedge \clk ) begin
        s375_val_n3 <= s374_val_n3;
    end
    always @(posedge \clk ) begin
        \s376_val  <= \s375_val ;
    end
    always @(posedge \clk ) begin
        s376_val_n1 <= s375_val_n1;
    end
    always @(posedge \clk ) begin
        s376_val_n2 <= s375_val_n2;
    end
    always @(posedge \clk ) begin
        s376_val_n3 <= s375_val_n3;
    end
    always @(posedge \clk ) begin
        \s377_val  <= \s376_val ;
    end
    always @(posedge \clk ) begin
        s377_val_n1 <= s376_val_n1;
    end
    always @(posedge \clk ) begin
        s377_val_n2 <= s376_val_n2;
    end
    always @(posedge \clk ) begin
        s377_val_n3 <= s376_val_n3;
    end
    always @(posedge \clk ) begin
        \s378_val  <= \s377_val ;
    end
    always @(posedge \clk ) begin
        s378_val_n1 <= s377_val_n1;
    end
    always @(posedge \clk ) begin
        s378_val_n2 <= s377_val_n2;
    end
    always @(posedge \clk ) begin
        s378_val_n3 <= s377_val_n3;
    end
    always @(posedge \clk ) begin
        \s379_val  <= \s378_val ;
    end
    always @(posedge \clk ) begin
        s379_val_n1 <= s378_val_n1;
    end
    always @(posedge \clk ) begin
        s379_val_n2 <= s378_val_n2;
    end
    always @(posedge \clk ) begin
        s379_val_n3 <= s378_val_n3;
    end
    always @(posedge \clk ) begin
        \s380_val  <= \s379_val ;
    end
    always @(posedge \clk ) begin
        s380_val_n1 <= s379_val_n1;
    end
    always @(posedge \clk ) begin
        s380_val_n2 <= s379_val_n2;
    end
    always @(posedge \clk ) begin
        s380_val_n3 <= s379_val_n3;
    end
    always @(posedge \clk ) begin
        \s381_val  <= \s380_val ;
    end
    always @(posedge \clk ) begin
        s381_val_n1 <= s380_val_n1;
    end
    always @(posedge \clk ) begin
        s381_val_n2 <= s380_val_n2;
    end
    always @(posedge \clk ) begin
        s381_val_n3 <= s380_val_n3;
    end
    always @(posedge \clk ) begin
        \s382_val  <= \s381_val ;
    end
    always @(posedge \clk ) begin
        s382_val_n1 <= s381_val_n1;
    end
    always @(posedge \clk ) begin
        s382_val_n2 <= s381_val_n2;
    end
    always @(posedge \clk ) begin
        s382_val_n3 <= s381_val_n3;
    end
    always @(posedge \clk ) begin
        \s383_val  <= \s382_val ;
    end
    always @(posedge \clk ) begin
        s383_val_n1 <= s382_val_n1;
    end
    always @(posedge \clk ) begin
        s383_val_n2 <= s382_val_n2;
    end
    always @(posedge \clk ) begin
        s383_val_n3 <= s382_val_n3;
    end
    always @(posedge \clk ) begin
        \s384_val  <= \s383_val ;
    end
    always @(posedge \clk ) begin
        s384_val_n1 <= s383_val_n1;
    end
    always @(posedge \clk ) begin
        s384_val_n2 <= s383_val_n2;
    end
    always @(posedge \clk ) begin
        s384_val_n3 <= s383_val_n3;
    end
    always @(posedge \clk ) begin
        \s385_val  <= \s384_val ;
    end
    always @(posedge \clk ) begin
        s385_val_n1 <= s384_val_n1;
    end
    always @(posedge \clk ) begin
        s385_val_n2 <= s384_val_n2;
    end
    always @(posedge \clk ) begin
        s385_val_n3 <= s384_val_n3;
    end
    always @(posedge \clk ) begin
        \s386_val  <= \s385_val ;
    end
    always @(posedge \clk ) begin
        s386_val_n1 <= s385_val_n1;
    end
    always @(posedge \clk ) begin
        s386_val_n2 <= s385_val_n2;
    end
    always @(posedge \clk ) begin
        s386_val_n3 <= s385_val_n3;
    end
    always @(posedge \clk ) begin
        \s387_val  <= \s386_val ;
    end
    always @(posedge \clk ) begin
        s387_val_n1 <= s386_val_n1;
    end
    always @(posedge \clk ) begin
        s387_val_n2 <= s386_val_n2;
    end
    always @(posedge \clk ) begin
        s387_val_n3 <= s386_val_n3;
    end
    always @(posedge \clk ) begin
        \s388_val  <= \s387_val ;
    end
    always @(posedge \clk ) begin
        s388_val_n1 <= s387_val_n1;
    end
    always @(posedge \clk ) begin
        s388_val_n2 <= s387_val_n2;
    end
    always @(posedge \clk ) begin
        s388_val_n3 <= s387_val_n3;
    end
    always @(posedge \clk ) begin
        \s389_val  <= \s388_val ;
    end
    always @(posedge \clk ) begin
        s389_val_n1 <= s388_val_n1;
    end
    always @(posedge \clk ) begin
        s389_val_n2 <= s388_val_n2;
    end
    always @(posedge \clk ) begin
        s389_val_n3 <= s388_val_n3;
    end
    always @(posedge \clk ) begin
        \s390_val  <= \s389_val ;
    end
    always @(posedge \clk ) begin
        s390_val_n1 <= s389_val_n1;
    end
    always @(posedge \clk ) begin
        s390_val_n2 <= s389_val_n2;
    end
    always @(posedge \clk ) begin
        s390_val_n3 <= s389_val_n3;
    end
    always @(posedge \clk ) begin
        \s391_val  <= \s390_val ;
    end
    always @(posedge \clk ) begin
        s391_val_n1 <= s390_val_n1;
    end
    always @(posedge \clk ) begin
        s391_val_n2 <= s390_val_n2;
    end
    always @(posedge \clk ) begin
        s391_val_n3 <= s390_val_n3;
    end
    always @(posedge \clk ) begin
        \s392_val  <= \s391_val ;
    end
    always @(posedge \clk ) begin
        s392_val_n1 <= s391_val_n1;
    end
    always @(posedge \clk ) begin
        s392_val_n2 <= s391_val_n2;
    end
    always @(posedge \clk ) begin
        s392_val_n3 <= s391_val_n3;
    end
    always @(posedge \clk ) begin
        \s393_val  <= \s392_val ;
    end
    always @(posedge \clk ) begin
        s393_val_n1 <= s392_val_n1;
    end
    always @(posedge \clk ) begin
        s393_val_n2 <= s392_val_n2;
    end
    always @(posedge \clk ) begin
        s393_val_n3 <= s392_val_n3;
    end
    always @(posedge \clk ) begin
        \s394_val  <= \s393_val ;
    end
    always @(posedge \clk ) begin
        s394_val_n1 <= s393_val_n1;
    end
    always @(posedge \clk ) begin
        s394_val_n2 <= s393_val_n2;
    end
    always @(posedge \clk ) begin
        s394_val_n3 <= s393_val_n3;
    end
    always @(posedge \clk ) begin
        \s395_val  <= \s394_val ;
    end
    always @(posedge \clk ) begin
        s395_val_n1 <= s394_val_n1;
    end
    always @(posedge \clk ) begin
        s395_val_n2 <= s394_val_n2;
    end
    always @(posedge \clk ) begin
        s395_val_n3 <= s394_val_n3;
    end
    always @(posedge \clk ) begin
        \s396_val  <= \s395_val ;
    end
    always @(posedge \clk ) begin
        s396_val_n1 <= s395_val_n1;
    end
    always @(posedge \clk ) begin
        s396_val_n2 <= s395_val_n2;
    end
    always @(posedge \clk ) begin
        s396_val_n3 <= s395_val_n3;
    end
    always @(posedge \clk ) begin
        \s397_val  <= \s396_val ;
    end
    always @(posedge \clk ) begin
        s397_val_n1 <= s396_val_n1;
    end
    always @(posedge \clk ) begin
        s397_val_n2 <= s396_val_n2;
    end
    always @(posedge \clk ) begin
        s397_val_n3 <= s396_val_n3;
    end
    always @(posedge \clk ) begin
        \s398_val  <= \s397_val ;
    end
    always @(posedge \clk ) begin
        s398_val_n1 <= s397_val_n1;
    end
    always @(posedge \clk ) begin
        s398_val_n2 <= s397_val_n2;
    end
    always @(posedge \clk ) begin
        s398_val_n3 <= s397_val_n3;
    end
    always @(posedge \clk ) begin
        \s399_val  <= \s398_val ;
    end
    always @(posedge \clk ) begin
        s399_val_n1 <= s398_val_n1;
    end
    always @(posedge \clk ) begin
        s399_val_n2 <= s398_val_n2;
    end
    always @(posedge \clk ) begin
        s399_val_n3 <= s398_val_n3;
    end
    always @(posedge \clk ) begin
        \s400_val  <= \s399_val ;
    end
    always @(posedge \clk ) begin
        s400_val_n1 <= s399_val_n1;
    end
    always @(posedge \clk ) begin
        s400_val_n2 <= s399_val_n2;
    end
    always @(posedge \clk ) begin
        s400_val_n3 <= s399_val_n3;
    end
    always @(posedge \clk ) begin
        \s401_val  <= \s400_val ;
    end
    always @(posedge \clk ) begin
        s401_val_n1 <= s400_val_n1;
    end
    always @(posedge \clk ) begin
        s401_val_n2 <= s400_val_n2;
    end
    always @(posedge \clk ) begin
        s401_val_n3 <= s400_val_n3;
    end
    always @(posedge \clk ) begin
        s401_val_n4 <= val_n4;
    end
    always @(posedge \clk ) begin
        \s402_val  <= \s401_val ;
    end
    always @(posedge \clk ) begin
        s402_val_n1 <= s401_val_n1;
    end
    always @(posedge \clk ) begin
        s402_val_n2 <= s401_val_n2;
    end
    always @(posedge \clk ) begin
        s402_val_n3 <= s401_val_n3;
    end
    always @(posedge \clk ) begin
        s402_val_n4 <= s401_val_n4;
    end
    always @(posedge \clk ) begin
        \s403_val  <= \s402_val ;
    end
    always @(posedge \clk ) begin
        s403_val_n1 <= s402_val_n1;
    end
    always @(posedge \clk ) begin
        s403_val_n2 <= s402_val_n2;
    end
    always @(posedge \clk ) begin
        s403_val_n3 <= s402_val_n3;
    end
    always @(posedge \clk ) begin
        s403_val_n4 <= s402_val_n4;
    end
    always @(posedge \clk ) begin
        \s404_val  <= \s403_val ;
    end
    always @(posedge \clk ) begin
        s404_val_n1 <= s403_val_n1;
    end
    always @(posedge \clk ) begin
        s404_val_n2 <= s403_val_n2;
    end
    always @(posedge \clk ) begin
        s404_val_n3 <= s403_val_n3;
    end
    always @(posedge \clk ) begin
        s404_val_n4 <= s403_val_n4;
    end
    always @(posedge \clk ) begin
        \s405_val  <= \s404_val ;
    end
    always @(posedge \clk ) begin
        s405_val_n1 <= s404_val_n1;
    end
    always @(posedge \clk ) begin
        s405_val_n2 <= s404_val_n2;
    end
    always @(posedge \clk ) begin
        s405_val_n3 <= s404_val_n3;
    end
    always @(posedge \clk ) begin
        s405_val_n4 <= s404_val_n4;
    end
    always @(posedge \clk ) begin
        \s406_val  <= \s405_val ;
    end
    always @(posedge \clk ) begin
        s406_val_n1 <= s405_val_n1;
    end
    always @(posedge \clk ) begin
        s406_val_n2 <= s405_val_n2;
    end
    always @(posedge \clk ) begin
        s406_val_n3 <= s405_val_n3;
    end
    always @(posedge \clk ) begin
        s406_val_n4 <= s405_val_n4;
    end
    always @(posedge \clk ) begin
        \s407_val  <= \s406_val ;
    end
    always @(posedge \clk ) begin
        s407_val_n1 <= s406_val_n1;
    end
    always @(posedge \clk ) begin
        s407_val_n2 <= s406_val_n2;
    end
    always @(posedge \clk ) begin
        s407_val_n3 <= s406_val_n3;
    end
    always @(posedge \clk ) begin
        s407_val_n4 <= s406_val_n4;
    end
    always @(posedge \clk ) begin
        \s408_val  <= \s407_val ;
    end
    always @(posedge \clk ) begin
        s408_val_n1 <= s407_val_n1;
    end
    always @(posedge \clk ) begin
        s408_val_n2 <= s407_val_n2;
    end
    always @(posedge \clk ) begin
        s408_val_n3 <= s407_val_n3;
    end
    always @(posedge \clk ) begin
        s408_val_n4 <= s407_val_n4;
    end
    always @(posedge \clk ) begin
        \s409_val  <= \s408_val ;
    end
    always @(posedge \clk ) begin
        s409_val_n1 <= s408_val_n1;
    end
    always @(posedge \clk ) begin
        s409_val_n2 <= s408_val_n2;
    end
    always @(posedge \clk ) begin
        s409_val_n3 <= s408_val_n3;
    end
    always @(posedge \clk ) begin
        s409_val_n4 <= s408_val_n4;
    end
    always @(posedge \clk ) begin
        \s410_val  <= \s409_val ;
    end
    always @(posedge \clk ) begin
        s410_val_n1 <= s409_val_n1;
    end
    always @(posedge \clk ) begin
        s410_val_n2 <= s409_val_n2;
    end
    always @(posedge \clk ) begin
        s410_val_n3 <= s409_val_n3;
    end
    always @(posedge \clk ) begin
        s410_val_n4 <= s409_val_n4;
    end
    always @(posedge \clk ) begin
        \s411_val  <= \s410_val ;
    end
    always @(posedge \clk ) begin
        s411_val_n1 <= s410_val_n1;
    end
    always @(posedge \clk ) begin
        s411_val_n2 <= s410_val_n2;
    end
    always @(posedge \clk ) begin
        s411_val_n3 <= s410_val_n3;
    end
    always @(posedge \clk ) begin
        s411_val_n4 <= s410_val_n4;
    end
    always @(posedge \clk ) begin
        \s412_val  <= \s411_val ;
    end
    always @(posedge \clk ) begin
        s412_val_n1 <= s411_val_n1;
    end
    always @(posedge \clk ) begin
        s412_val_n2 <= s411_val_n2;
    end
    always @(posedge \clk ) begin
        s412_val_n3 <= s411_val_n3;
    end
    always @(posedge \clk ) begin
        s412_val_n4 <= s411_val_n4;
    end
    always @(posedge \clk ) begin
        \s413_val  <= \s412_val ;
    end
    always @(posedge \clk ) begin
        s413_val_n1 <= s412_val_n1;
    end
    always @(posedge \clk ) begin
        s413_val_n2 <= s412_val_n2;
    end
    always @(posedge \clk ) begin
        s413_val_n3 <= s412_val_n3;
    end
    always @(posedge \clk ) begin
        s413_val_n4 <= s412_val_n4;
    end
    always @(posedge \clk ) begin
        \s414_val  <= \s413_val ;
    end
    always @(posedge \clk ) begin
        s414_val_n1 <= s413_val_n1;
    end
    always @(posedge \clk ) begin
        s414_val_n2 <= s413_val_n2;
    end
    always @(posedge \clk ) begin
        s414_val_n3 <= s413_val_n3;
    end
    always @(posedge \clk ) begin
        s414_val_n4 <= s413_val_n4;
    end
    always @(posedge \clk ) begin
        \s415_val  <= \s414_val ;
    end
    always @(posedge \clk ) begin
        s415_val_n1 <= s414_val_n1;
    end
    always @(posedge \clk ) begin
        s415_val_n2 <= s414_val_n2;
    end
    always @(posedge \clk ) begin
        s415_val_n3 <= s414_val_n3;
    end
    always @(posedge \clk ) begin
        s415_val_n4 <= s414_val_n4;
    end
    always @(posedge \clk ) begin
        \s416_val  <= \s415_val ;
    end
    always @(posedge \clk ) begin
        s416_val_n1 <= s415_val_n1;
    end
    always @(posedge \clk ) begin
        s416_val_n2 <= s415_val_n2;
    end
    always @(posedge \clk ) begin
        s416_val_n3 <= s415_val_n3;
    end
    always @(posedge \clk ) begin
        s416_val_n4 <= s415_val_n4;
    end
    always @(posedge \clk ) begin
        \s417_val  <= \s416_val ;
    end
    always @(posedge \clk ) begin
        s417_val_n1 <= s416_val_n1;
    end
    always @(posedge \clk ) begin
        s417_val_n2 <= s416_val_n2;
    end
    always @(posedge \clk ) begin
        s417_val_n3 <= s416_val_n3;
    end
    always @(posedge \clk ) begin
        s417_val_n4 <= s416_val_n4;
    end
    always @(posedge \clk ) begin
        \s418_val  <= \s417_val ;
    end
    always @(posedge \clk ) begin
        s418_val_n1 <= s417_val_n1;
    end
    always @(posedge \clk ) begin
        s418_val_n2 <= s417_val_n2;
    end
    always @(posedge \clk ) begin
        s418_val_n3 <= s417_val_n3;
    end
    always @(posedge \clk ) begin
        s418_val_n4 <= s417_val_n4;
    end
    always @(posedge \clk ) begin
        \s419_val  <= \s418_val ;
    end
    always @(posedge \clk ) begin
        s419_val_n1 <= s418_val_n1;
    end
    always @(posedge \clk ) begin
        s419_val_n2 <= s418_val_n2;
    end
    always @(posedge \clk ) begin
        s419_val_n3 <= s418_val_n3;
    end
    always @(posedge \clk ) begin
        s419_val_n4 <= s418_val_n4;
    end
    always @(posedge \clk ) begin
        \s420_val  <= \s419_val ;
    end
    always @(posedge \clk ) begin
        s420_val_n1 <= s419_val_n1;
    end
    always @(posedge \clk ) begin
        s420_val_n2 <= s419_val_n2;
    end
    always @(posedge \clk ) begin
        s420_val_n3 <= s419_val_n3;
    end
    always @(posedge \clk ) begin
        s420_val_n4 <= s419_val_n4;
    end
    always @(posedge \clk ) begin
        \s421_val  <= \s420_val ;
    end
    always @(posedge \clk ) begin
        s421_val_n1 <= s420_val_n1;
    end
    always @(posedge \clk ) begin
        s421_val_n2 <= s420_val_n2;
    end
    always @(posedge \clk ) begin
        s421_val_n3 <= s420_val_n3;
    end
    always @(posedge \clk ) begin
        s421_val_n4 <= s420_val_n4;
    end
    always @(posedge \clk ) begin
        \s422_val  <= \s421_val ;
    end
    always @(posedge \clk ) begin
        s422_val_n1 <= s421_val_n1;
    end
    always @(posedge \clk ) begin
        s422_val_n2 <= s421_val_n2;
    end
    always @(posedge \clk ) begin
        s422_val_n3 <= s421_val_n3;
    end
    always @(posedge \clk ) begin
        s422_val_n4 <= s421_val_n4;
    end
    always @(posedge \clk ) begin
        \s423_val  <= \s422_val ;
    end
    always @(posedge \clk ) begin
        s423_val_n1 <= s422_val_n1;
    end
    always @(posedge \clk ) begin
        s423_val_n2 <= s422_val_n2;
    end
    always @(posedge \clk ) begin
        s423_val_n3 <= s422_val_n3;
    end
    always @(posedge \clk ) begin
        s423_val_n4 <= s422_val_n4;
    end
    always @(posedge \clk ) begin
        \s424_val  <= \s423_val ;
    end
    always @(posedge \clk ) begin
        s424_val_n1 <= s423_val_n1;
    end
    always @(posedge \clk ) begin
        s424_val_n2 <= s423_val_n2;
    end
    always @(posedge \clk ) begin
        s424_val_n3 <= s423_val_n3;
    end
    always @(posedge \clk ) begin
        s424_val_n4 <= s423_val_n4;
    end
    always @(posedge \clk ) begin
        \s425_val  <= \s424_val ;
    end
    always @(posedge \clk ) begin
        s425_val_n1 <= s424_val_n1;
    end
    always @(posedge \clk ) begin
        s425_val_n2 <= s424_val_n2;
    end
    always @(posedge \clk ) begin
        s425_val_n3 <= s424_val_n3;
    end
    always @(posedge \clk ) begin
        s425_val_n4 <= s424_val_n4;
    end
    always @(posedge \clk ) begin
        \s426_val  <= \s425_val ;
    end
    always @(posedge \clk ) begin
        s426_val_n1 <= s425_val_n1;
    end
    always @(posedge \clk ) begin
        s426_val_n2 <= s425_val_n2;
    end
    always @(posedge \clk ) begin
        s426_val_n3 <= s425_val_n3;
    end
    always @(posedge \clk ) begin
        s426_val_n4 <= s425_val_n4;
    end
    always @(posedge \clk ) begin
        \s427_val  <= \s426_val ;
    end
    always @(posedge \clk ) begin
        s427_val_n1 <= s426_val_n1;
    end
    always @(posedge \clk ) begin
        s427_val_n2 <= s426_val_n2;
    end
    always @(posedge \clk ) begin
        s427_val_n3 <= s426_val_n3;
    end
    always @(posedge \clk ) begin
        s427_val_n4 <= s426_val_n4;
    end
    always @(posedge \clk ) begin
        \s428_val  <= \s427_val ;
    end
    always @(posedge \clk ) begin
        s428_val_n1 <= s427_val_n1;
    end
    always @(posedge \clk ) begin
        s428_val_n2 <= s427_val_n2;
    end
    always @(posedge \clk ) begin
        s428_val_n3 <= s427_val_n3;
    end
    always @(posedge \clk ) begin
        s428_val_n4 <= s427_val_n4;
    end
    always @(posedge \clk ) begin
        \s429_val  <= \s428_val ;
    end
    always @(posedge \clk ) begin
        s429_val_n1 <= s428_val_n1;
    end
    always @(posedge \clk ) begin
        s429_val_n2 <= s428_val_n2;
    end
    always @(posedge \clk ) begin
        s429_val_n3 <= s428_val_n3;
    end
    always @(posedge \clk ) begin
        s429_val_n4 <= s428_val_n4;
    end
    always @(posedge \clk ) begin
        \s430_val  <= \s429_val ;
    end
    always @(posedge \clk ) begin
        s430_val_n1 <= s429_val_n1;
    end
    always @(posedge \clk ) begin
        s430_val_n2 <= s429_val_n2;
    end
    always @(posedge \clk ) begin
        s430_val_n3 <= s429_val_n3;
    end
    always @(posedge \clk ) begin
        s430_val_n4 <= s429_val_n4;
    end
    always @(posedge \clk ) begin
        \s431_val  <= \s430_val ;
    end
    always @(posedge \clk ) begin
        s431_val_n1 <= s430_val_n1;
    end
    always @(posedge \clk ) begin
        s431_val_n2 <= s430_val_n2;
    end
    always @(posedge \clk ) begin
        s431_val_n3 <= s430_val_n3;
    end
    always @(posedge \clk ) begin
        s431_val_n4 <= s430_val_n4;
    end
    always @(posedge \clk ) begin
        \s432_val  <= \s431_val ;
    end
    always @(posedge \clk ) begin
        s432_val_n1 <= s431_val_n1;
    end
    always @(posedge \clk ) begin
        s432_val_n2 <= s431_val_n2;
    end
    always @(posedge \clk ) begin
        s432_val_n3 <= s431_val_n3;
    end
    always @(posedge \clk ) begin
        s432_val_n4 <= s431_val_n4;
    end
    always @(posedge \clk ) begin
        \s433_val  <= \s432_val ;
    end
    always @(posedge \clk ) begin
        s433_val_n1 <= s432_val_n1;
    end
    always @(posedge \clk ) begin
        s433_val_n2 <= s432_val_n2;
    end
    always @(posedge \clk ) begin
        s433_val_n3 <= s432_val_n3;
    end
    always @(posedge \clk ) begin
        s433_val_n4 <= s432_val_n4;
    end
    always @(posedge \clk ) begin
        \s434_val  <= \s433_val ;
    end
    always @(posedge \clk ) begin
        s434_val_n1 <= s433_val_n1;
    end
    always @(posedge \clk ) begin
        s434_val_n2 <= s433_val_n2;
    end
    always @(posedge \clk ) begin
        s434_val_n3 <= s433_val_n3;
    end
    always @(posedge \clk ) begin
        s434_val_n4 <= s433_val_n4;
    end
    always @(posedge \clk ) begin
        \s435_val  <= \s434_val ;
    end
    always @(posedge \clk ) begin
        s435_val_n1 <= s434_val_n1;
    end
    always @(posedge \clk ) begin
        s435_val_n2 <= s434_val_n2;
    end
    always @(posedge \clk ) begin
        s435_val_n3 <= s434_val_n3;
    end
    always @(posedge \clk ) begin
        s435_val_n4 <= s434_val_n4;
    end
    always @(posedge \clk ) begin
        \s436_val  <= \s435_val ;
    end
    always @(posedge \clk ) begin
        s436_val_n1 <= s435_val_n1;
    end
    always @(posedge \clk ) begin
        s436_val_n2 <= s435_val_n2;
    end
    always @(posedge \clk ) begin
        s436_val_n3 <= s435_val_n3;
    end
    always @(posedge \clk ) begin
        s436_val_n4 <= s435_val_n4;
    end
    always @(posedge \clk ) begin
        \s437_val  <= \s436_val ;
    end
    always @(posedge \clk ) begin
        s437_val_n1 <= s436_val_n1;
    end
    always @(posedge \clk ) begin
        s437_val_n2 <= s436_val_n2;
    end
    always @(posedge \clk ) begin
        s437_val_n3 <= s436_val_n3;
    end
    always @(posedge \clk ) begin
        s437_val_n4 <= s436_val_n4;
    end
    always @(posedge \clk ) begin
        \s438_val  <= \s437_val ;
    end
    always @(posedge \clk ) begin
        s438_val_n1 <= s437_val_n1;
    end
    always @(posedge \clk ) begin
        s438_val_n2 <= s437_val_n2;
    end
    always @(posedge \clk ) begin
        s438_val_n3 <= s437_val_n3;
    end
    always @(posedge \clk ) begin
        s438_val_n4 <= s437_val_n4;
    end
    always @(posedge \clk ) begin
        \s439_val  <= \s438_val ;
    end
    always @(posedge \clk ) begin
        s439_val_n1 <= s438_val_n1;
    end
    always @(posedge \clk ) begin
        s439_val_n2 <= s438_val_n2;
    end
    always @(posedge \clk ) begin
        s439_val_n3 <= s438_val_n3;
    end
    always @(posedge \clk ) begin
        s439_val_n4 <= s438_val_n4;
    end
    always @(posedge \clk ) begin
        \s440_val  <= \s439_val ;
    end
    always @(posedge \clk ) begin
        s440_val_n1 <= s439_val_n1;
    end
    always @(posedge \clk ) begin
        s440_val_n2 <= s439_val_n2;
    end
    always @(posedge \clk ) begin
        s440_val_n3 <= s439_val_n3;
    end
    always @(posedge \clk ) begin
        s440_val_n4 <= s439_val_n4;
    end
    always @(posedge \clk ) begin
        \s441_val  <= \s440_val ;
    end
    always @(posedge \clk ) begin
        s441_val_n1 <= s440_val_n1;
    end
    always @(posedge \clk ) begin
        s441_val_n2 <= s440_val_n2;
    end
    always @(posedge \clk ) begin
        s441_val_n3 <= s440_val_n3;
    end
    always @(posedge \clk ) begin
        s441_val_n4 <= s440_val_n4;
    end
    always @(posedge \clk ) begin
        \s442_val  <= \s441_val ;
    end
    always @(posedge \clk ) begin
        s442_val_n1 <= s441_val_n1;
    end
    always @(posedge \clk ) begin
        s442_val_n2 <= s441_val_n2;
    end
    always @(posedge \clk ) begin
        s442_val_n3 <= s441_val_n3;
    end
    always @(posedge \clk ) begin
        s442_val_n4 <= s441_val_n4;
    end
    always @(posedge \clk ) begin
        \s443_val  <= \s442_val ;
    end
    always @(posedge \clk ) begin
        s443_val_n1 <= s442_val_n1;
    end
    always @(posedge \clk ) begin
        s443_val_n2 <= s442_val_n2;
    end
    always @(posedge \clk ) begin
        s443_val_n3 <= s442_val_n3;
    end
    always @(posedge \clk ) begin
        s443_val_n4 <= s442_val_n4;
    end
    always @(posedge \clk ) begin
        \s444_val  <= \s443_val ;
    end
    always @(posedge \clk ) begin
        s444_val_n1 <= s443_val_n1;
    end
    always @(posedge \clk ) begin
        s444_val_n2 <= s443_val_n2;
    end
    always @(posedge \clk ) begin
        s444_val_n3 <= s443_val_n3;
    end
    always @(posedge \clk ) begin
        s444_val_n4 <= s443_val_n4;
    end
    always @(posedge \clk ) begin
        \s445_val  <= \s444_val ;
    end
    always @(posedge \clk ) begin
        s445_val_n1 <= s444_val_n1;
    end
    always @(posedge \clk ) begin
        s445_val_n2 <= s444_val_n2;
    end
    always @(posedge \clk ) begin
        s445_val_n3 <= s444_val_n3;
    end
    always @(posedge \clk ) begin
        s445_val_n4 <= s444_val_n4;
    end
    always @(posedge \clk ) begin
        \s446_val  <= \s445_val ;
    end
    always @(posedge \clk ) begin
        s446_val_n1 <= s445_val_n1;
    end
    always @(posedge \clk ) begin
        s446_val_n2 <= s445_val_n2;
    end
    always @(posedge \clk ) begin
        s446_val_n3 <= s445_val_n3;
    end
    always @(posedge \clk ) begin
        s446_val_n4 <= s445_val_n4;
    end
    always @(posedge \clk ) begin
        \s447_val  <= \s446_val ;
    end
    always @(posedge \clk ) begin
        s447_val_n1 <= s446_val_n1;
    end
    always @(posedge \clk ) begin
        s447_val_n2 <= s446_val_n2;
    end
    always @(posedge \clk ) begin
        s447_val_n3 <= s446_val_n3;
    end
    always @(posedge \clk ) begin
        s447_val_n4 <= s446_val_n4;
    end
    always @(posedge \clk ) begin
        \s448_val  <= \s447_val ;
    end
    always @(posedge \clk ) begin
        s448_val_n1 <= s447_val_n1;
    end
    always @(posedge \clk ) begin
        s448_val_n2 <= s447_val_n2;
    end
    always @(posedge \clk ) begin
        s448_val_n3 <= s447_val_n3;
    end
    always @(posedge \clk ) begin
        s448_val_n4 <= s447_val_n4;
    end
    always @(posedge \clk ) begin
        \s449_val  <= \s448_val ;
    end
    always @(posedge \clk ) begin
        s449_val_n1 <= s448_val_n1;
    end
    always @(posedge \clk ) begin
        s449_val_n2 <= s448_val_n2;
    end
    always @(posedge \clk ) begin
        s449_val_n3 <= s448_val_n3;
    end
    always @(posedge \clk ) begin
        s449_val_n4 <= s448_val_n4;
    end
    always @(posedge \clk ) begin
        \s450_val  <= \s449_val ;
    end
    always @(posedge \clk ) begin
        s450_val_n1 <= s449_val_n1;
    end
    always @(posedge \clk ) begin
        s450_val_n2 <= s449_val_n2;
    end
    always @(posedge \clk ) begin
        s450_val_n3 <= s449_val_n3;
    end
    always @(posedge \clk ) begin
        s450_val_n4 <= s449_val_n4;
    end
    always @(posedge \clk ) begin
        \s451_val  <= \s450_val ;
    end
    always @(posedge \clk ) begin
        s451_val_n1 <= s450_val_n1;
    end
    always @(posedge \clk ) begin
        s451_val_n2 <= s450_val_n2;
    end
    always @(posedge \clk ) begin
        s451_val_n3 <= s450_val_n3;
    end
    always @(posedge \clk ) begin
        s451_val_n4 <= s450_val_n4;
    end
    always @(posedge \clk ) begin
        \s452_val  <= \s451_val ;
    end
    always @(posedge \clk ) begin
        s452_val_n1 <= s451_val_n1;
    end
    always @(posedge \clk ) begin
        s452_val_n2 <= s451_val_n2;
    end
    always @(posedge \clk ) begin
        s452_val_n3 <= s451_val_n3;
    end
    always @(posedge \clk ) begin
        s452_val_n4 <= s451_val_n4;
    end
    always @(posedge \clk ) begin
        \s453_val  <= \s452_val ;
    end
    always @(posedge \clk ) begin
        s453_val_n1 <= s452_val_n1;
    end
    always @(posedge \clk ) begin
        s453_val_n2 <= s452_val_n2;
    end
    always @(posedge \clk ) begin
        s453_val_n3 <= s452_val_n3;
    end
    always @(posedge \clk ) begin
        s453_val_n4 <= s452_val_n4;
    end
    always @(posedge \clk ) begin
        \s454_val  <= \s453_val ;
    end
    always @(posedge \clk ) begin
        s454_val_n1 <= s453_val_n1;
    end
    always @(posedge \clk ) begin
        s454_val_n2 <= s453_val_n2;
    end
    always @(posedge \clk ) begin
        s454_val_n3 <= s453_val_n3;
    end
    always @(posedge \clk ) begin
        s454_val_n4 <= s453_val_n4;
    end
    always @(posedge \clk ) begin
        \s455_val  <= \s454_val ;
    end
    always @(posedge \clk ) begin
        s455_val_n1 <= s454_val_n1;
    end
    always @(posedge \clk ) begin
        s455_val_n2 <= s454_val_n2;
    end
    always @(posedge \clk ) begin
        s455_val_n3 <= s454_val_n3;
    end
    always @(posedge \clk ) begin
        s455_val_n4 <= s454_val_n4;
    end
    always @(posedge \clk ) begin
        \s456_val  <= \s455_val ;
    end
    always @(posedge \clk ) begin
        s456_val_n1 <= s455_val_n1;
    end
    always @(posedge \clk ) begin
        s456_val_n2 <= s455_val_n2;
    end
    always @(posedge \clk ) begin
        s456_val_n3 <= s455_val_n3;
    end
    always @(posedge \clk ) begin
        s456_val_n4 <= s455_val_n4;
    end
    always @(posedge \clk ) begin
        \s457_val  <= \s456_val ;
    end
    always @(posedge \clk ) begin
        s457_val_n1 <= s456_val_n1;
    end
    always @(posedge \clk ) begin
        s457_val_n2 <= s456_val_n2;
    end
    always @(posedge \clk ) begin
        s457_val_n3 <= s456_val_n3;
    end
    always @(posedge \clk ) begin
        s457_val_n4 <= s456_val_n4;
    end
    always @(posedge \clk ) begin
        \s458_val  <= \s457_val ;
    end
    always @(posedge \clk ) begin
        s458_val_n1 <= s457_val_n1;
    end
    always @(posedge \clk ) begin
        s458_val_n2 <= s457_val_n2;
    end
    always @(posedge \clk ) begin
        s458_val_n3 <= s457_val_n3;
    end
    always @(posedge \clk ) begin
        s458_val_n4 <= s457_val_n4;
    end
    always @(posedge \clk ) begin
        \s459_val  <= \s458_val ;
    end
    always @(posedge \clk ) begin
        s459_val_n1 <= s458_val_n1;
    end
    always @(posedge \clk ) begin
        s459_val_n2 <= s458_val_n2;
    end
    always @(posedge \clk ) begin
        s459_val_n3 <= s458_val_n3;
    end
    always @(posedge \clk ) begin
        s459_val_n4 <= s458_val_n4;
    end
    always @(posedge \clk ) begin
        \s460_val  <= \s459_val ;
    end
    always @(posedge \clk ) begin
        s460_val_n1 <= s459_val_n1;
    end
    always @(posedge \clk ) begin
        s460_val_n2 <= s459_val_n2;
    end
    always @(posedge \clk ) begin
        s460_val_n3 <= s459_val_n3;
    end
    always @(posedge \clk ) begin
        s460_val_n4 <= s459_val_n4;
    end
    always @(posedge \clk ) begin
        \s461_val  <= \s460_val ;
    end
    always @(posedge \clk ) begin
        s461_val_n1 <= s460_val_n1;
    end
    always @(posedge \clk ) begin
        s461_val_n2 <= s460_val_n2;
    end
    always @(posedge \clk ) begin
        s461_val_n3 <= s460_val_n3;
    end
    always @(posedge \clk ) begin
        s461_val_n4 <= s460_val_n4;
    end
    always @(posedge \clk ) begin
        \s462_val  <= \s461_val ;
    end
    always @(posedge \clk ) begin
        s462_val_n1 <= s461_val_n1;
    end
    always @(posedge \clk ) begin
        s462_val_n2 <= s461_val_n2;
    end
    always @(posedge \clk ) begin
        s462_val_n3 <= s461_val_n3;
    end
    always @(posedge \clk ) begin
        s462_val_n4 <= s461_val_n4;
    end
    always @(posedge \clk ) begin
        \s463_val  <= \s462_val ;
    end
    always @(posedge \clk ) begin
        s463_val_n1 <= s462_val_n1;
    end
    always @(posedge \clk ) begin
        s463_val_n2 <= s462_val_n2;
    end
    always @(posedge \clk ) begin
        s463_val_n3 <= s462_val_n3;
    end
    always @(posedge \clk ) begin
        s463_val_n4 <= s462_val_n4;
    end
    always @(posedge \clk ) begin
        \s464_val  <= \s463_val ;
    end
    always @(posedge \clk ) begin
        s464_val_n1 <= s463_val_n1;
    end
    always @(posedge \clk ) begin
        s464_val_n2 <= s463_val_n2;
    end
    always @(posedge \clk ) begin
        s464_val_n3 <= s463_val_n3;
    end
    always @(posedge \clk ) begin
        s464_val_n4 <= s463_val_n4;
    end
    always @(posedge \clk ) begin
        \s465_val  <= \s464_val ;
    end
    always @(posedge \clk ) begin
        s465_val_n1 <= s464_val_n1;
    end
    always @(posedge \clk ) begin
        s465_val_n2 <= s464_val_n2;
    end
    always @(posedge \clk ) begin
        s465_val_n3 <= s464_val_n3;
    end
    always @(posedge \clk ) begin
        s465_val_n4 <= s464_val_n4;
    end
    always @(posedge \clk ) begin
        \s466_val  <= \s465_val ;
    end
    always @(posedge \clk ) begin
        s466_val_n1 <= s465_val_n1;
    end
    always @(posedge \clk ) begin
        s466_val_n2 <= s465_val_n2;
    end
    always @(posedge \clk ) begin
        s466_val_n3 <= s465_val_n3;
    end
    always @(posedge \clk ) begin
        s466_val_n4 <= s465_val_n4;
    end
    always @(posedge \clk ) begin
        \s467_val  <= \s466_val ;
    end
    always @(posedge \clk ) begin
        s467_val_n1 <= s466_val_n1;
    end
    always @(posedge \clk ) begin
        s467_val_n2 <= s466_val_n2;
    end
    always @(posedge \clk ) begin
        s467_val_n3 <= s466_val_n3;
    end
    always @(posedge \clk ) begin
        s467_val_n4 <= s466_val_n4;
    end
    always @(posedge \clk ) begin
        \s468_val  <= \s467_val ;
    end
    always @(posedge \clk ) begin
        s468_val_n1 <= s467_val_n1;
    end
    always @(posedge \clk ) begin
        s468_val_n2 <= s467_val_n2;
    end
    always @(posedge \clk ) begin
        s468_val_n3 <= s467_val_n3;
    end
    always @(posedge \clk ) begin
        s468_val_n4 <= s467_val_n4;
    end
    always @(posedge \clk ) begin
        \s469_val  <= \s468_val ;
    end
    always @(posedge \clk ) begin
        s469_val_n1 <= s468_val_n1;
    end
    always @(posedge \clk ) begin
        s469_val_n2 <= s468_val_n2;
    end
    always @(posedge \clk ) begin
        s469_val_n3 <= s468_val_n3;
    end
    always @(posedge \clk ) begin
        s469_val_n4 <= s468_val_n4;
    end
    always @(posedge \clk ) begin
        \s470_val  <= \s469_val ;
    end
    always @(posedge \clk ) begin
        s470_val_n1 <= s469_val_n1;
    end
    always @(posedge \clk ) begin
        s470_val_n2 <= s469_val_n2;
    end
    always @(posedge \clk ) begin
        s470_val_n3 <= s469_val_n3;
    end
    always @(posedge \clk ) begin
        s470_val_n4 <= s469_val_n4;
    end
    always @(posedge \clk ) begin
        \s471_val  <= \s470_val ;
    end
    always @(posedge \clk ) begin
        s471_val_n1 <= s470_val_n1;
    end
    always @(posedge \clk ) begin
        s471_val_n2 <= s470_val_n2;
    end
    always @(posedge \clk ) begin
        s471_val_n3 <= s470_val_n3;
    end
    always @(posedge \clk ) begin
        s471_val_n4 <= s470_val_n4;
    end
    always @(posedge \clk ) begin
        \s472_val  <= \s471_val ;
    end
    always @(posedge \clk ) begin
        s472_val_n1 <= s471_val_n1;
    end
    always @(posedge \clk ) begin
        s472_val_n2 <= s471_val_n2;
    end
    always @(posedge \clk ) begin
        s472_val_n3 <= s471_val_n3;
    end
    always @(posedge \clk ) begin
        s472_val_n4 <= s471_val_n4;
    end
    always @(posedge \clk ) begin
        \s473_val  <= \s472_val ;
    end
    always @(posedge \clk ) begin
        s473_val_n1 <= s472_val_n1;
    end
    always @(posedge \clk ) begin
        s473_val_n2 <= s472_val_n2;
    end
    always @(posedge \clk ) begin
        s473_val_n3 <= s472_val_n3;
    end
    always @(posedge \clk ) begin
        s473_val_n4 <= s472_val_n4;
    end
    always @(posedge \clk ) begin
        \s474_val  <= \s473_val ;
    end
    always @(posedge \clk ) begin
        s474_val_n1 <= s473_val_n1;
    end
    always @(posedge \clk ) begin
        s474_val_n2 <= s473_val_n2;
    end
    always @(posedge \clk ) begin
        s474_val_n3 <= s473_val_n3;
    end
    always @(posedge \clk ) begin
        s474_val_n4 <= s473_val_n4;
    end
    always @(posedge \clk ) begin
        \s475_val  <= \s474_val ;
    end
    always @(posedge \clk ) begin
        s475_val_n1 <= s474_val_n1;
    end
    always @(posedge \clk ) begin
        s475_val_n2 <= s474_val_n2;
    end
    always @(posedge \clk ) begin
        s475_val_n3 <= s474_val_n3;
    end
    always @(posedge \clk ) begin
        s475_val_n4 <= s474_val_n4;
    end
    always @(posedge \clk ) begin
        \s476_val  <= \s475_val ;
    end
    always @(posedge \clk ) begin
        s476_val_n1 <= s475_val_n1;
    end
    always @(posedge \clk ) begin
        s476_val_n2 <= s475_val_n2;
    end
    always @(posedge \clk ) begin
        s476_val_n3 <= s475_val_n3;
    end
    always @(posedge \clk ) begin
        s476_val_n4 <= s475_val_n4;
    end
    always @(posedge \clk ) begin
        \s477_val  <= \s476_val ;
    end
    always @(posedge \clk ) begin
        s477_val_n1 <= s476_val_n1;
    end
    always @(posedge \clk ) begin
        s477_val_n2 <= s476_val_n2;
    end
    always @(posedge \clk ) begin
        s477_val_n3 <= s476_val_n3;
    end
    always @(posedge \clk ) begin
        s477_val_n4 <= s476_val_n4;
    end
    always @(posedge \clk ) begin
        \s478_val  <= \s477_val ;
    end
    always @(posedge \clk ) begin
        s478_val_n1 <= s477_val_n1;
    end
    always @(posedge \clk ) begin
        s478_val_n2 <= s477_val_n2;
    end
    always @(posedge \clk ) begin
        s478_val_n3 <= s477_val_n3;
    end
    always @(posedge \clk ) begin
        s478_val_n4 <= s477_val_n4;
    end
    always @(posedge \clk ) begin
        \s479_val  <= \s478_val ;
    end
    always @(posedge \clk ) begin
        s479_val_n1 <= s478_val_n1;
    end
    always @(posedge \clk ) begin
        s479_val_n2 <= s478_val_n2;
    end
    always @(posedge \clk ) begin
        s479_val_n3 <= s478_val_n3;
    end
    always @(posedge \clk ) begin
        s479_val_n4 <= s478_val_n4;
    end
    always @(posedge \clk ) begin
        \s480_val  <= \s479_val ;
    end
    always @(posedge \clk ) begin
        s480_val_n1 <= s479_val_n1;
    end
    always @(posedge \clk ) begin
        s480_val_n2 <= s479_val_n2;
    end
    always @(posedge \clk ) begin
        s480_val_n3 <= s479_val_n3;
    end
    always @(posedge \clk ) begin
        s480_val_n4 <= s479_val_n4;
    end
    always @(posedge \clk ) begin
        \s481_val  <= \s480_val ;
    end
    always @(posedge \clk ) begin
        s481_val_n1 <= s480_val_n1;
    end
    always @(posedge \clk ) begin
        s481_val_n2 <= s480_val_n2;
    end
    always @(posedge \clk ) begin
        s481_val_n3 <= s480_val_n3;
    end
    always @(posedge \clk ) begin
        s481_val_n4 <= s480_val_n4;
    end
    always @(posedge \clk ) begin
        \s482_val  <= \s481_val ;
    end
    always @(posedge \clk ) begin
        s482_val_n1 <= s481_val_n1;
    end
    always @(posedge \clk ) begin
        s482_val_n2 <= s481_val_n2;
    end
    always @(posedge \clk ) begin
        s482_val_n3 <= s481_val_n3;
    end
    always @(posedge \clk ) begin
        s482_val_n4 <= s481_val_n4;
    end
    always @(posedge \clk ) begin
        \s483_val  <= \s482_val ;
    end
    always @(posedge \clk ) begin
        s483_val_n1 <= s482_val_n1;
    end
    always @(posedge \clk ) begin
        s483_val_n2 <= s482_val_n2;
    end
    always @(posedge \clk ) begin
        s483_val_n3 <= s482_val_n3;
    end
    always @(posedge \clk ) begin
        s483_val_n4 <= s482_val_n4;
    end
    always @(posedge \clk ) begin
        \s484_val  <= \s483_val ;
    end
    always @(posedge \clk ) begin
        s484_val_n1 <= s483_val_n1;
    end
    always @(posedge \clk ) begin
        s484_val_n2 <= s483_val_n2;
    end
    always @(posedge \clk ) begin
        s484_val_n3 <= s483_val_n3;
    end
    always @(posedge \clk ) begin
        s484_val_n4 <= s483_val_n4;
    end
    always @(posedge \clk ) begin
        \s485_val  <= \s484_val ;
    end
    always @(posedge \clk ) begin
        s485_val_n1 <= s484_val_n1;
    end
    always @(posedge \clk ) begin
        s485_val_n2 <= s484_val_n2;
    end
    always @(posedge \clk ) begin
        s485_val_n3 <= s484_val_n3;
    end
    always @(posedge \clk ) begin
        s485_val_n4 <= s484_val_n4;
    end
    always @(posedge \clk ) begin
        \s486_val  <= \s485_val ;
    end
    always @(posedge \clk ) begin
        s486_val_n1 <= s485_val_n1;
    end
    always @(posedge \clk ) begin
        s486_val_n2 <= s485_val_n2;
    end
    always @(posedge \clk ) begin
        s486_val_n3 <= s485_val_n3;
    end
    always @(posedge \clk ) begin
        s486_val_n4 <= s485_val_n4;
    end
    always @(posedge \clk ) begin
        \s487_val  <= \s486_val ;
    end
    always @(posedge \clk ) begin
        s487_val_n1 <= s486_val_n1;
    end
    always @(posedge \clk ) begin
        s487_val_n2 <= s486_val_n2;
    end
    always @(posedge \clk ) begin
        s487_val_n3 <= s486_val_n3;
    end
    always @(posedge \clk ) begin
        s487_val_n4 <= s486_val_n4;
    end
    always @(posedge \clk ) begin
        \s488_val  <= \s487_val ;
    end
    always @(posedge \clk ) begin
        s488_val_n1 <= s487_val_n1;
    end
    always @(posedge \clk ) begin
        s488_val_n2 <= s487_val_n2;
    end
    always @(posedge \clk ) begin
        s488_val_n3 <= s487_val_n3;
    end
    always @(posedge \clk ) begin
        s488_val_n4 <= s487_val_n4;
    end
    always @(posedge \clk ) begin
        \s489_val  <= \s488_val ;
    end
    always @(posedge \clk ) begin
        s489_val_n1 <= s488_val_n1;
    end
    always @(posedge \clk ) begin
        s489_val_n2 <= s488_val_n2;
    end
    always @(posedge \clk ) begin
        s489_val_n3 <= s488_val_n3;
    end
    always @(posedge \clk ) begin
        s489_val_n4 <= s488_val_n4;
    end
    always @(posedge \clk ) begin
        \s490_val  <= \s489_val ;
    end
    always @(posedge \clk ) begin
        s490_val_n1 <= s489_val_n1;
    end
    always @(posedge \clk ) begin
        s490_val_n2 <= s489_val_n2;
    end
    always @(posedge \clk ) begin
        s490_val_n3 <= s489_val_n3;
    end
    always @(posedge \clk ) begin
        s490_val_n4 <= s489_val_n4;
    end
    always @(posedge \clk ) begin
        \s491_val  <= \s490_val ;
    end
    always @(posedge \clk ) begin
        s491_val_n1 <= s490_val_n1;
    end
    always @(posedge \clk ) begin
        s491_val_n2 <= s490_val_n2;
    end
    always @(posedge \clk ) begin
        s491_val_n3 <= s490_val_n3;
    end
    always @(posedge \clk ) begin
        s491_val_n4 <= s490_val_n4;
    end
    always @(posedge \clk ) begin
        \s492_val  <= \s491_val ;
    end
    always @(posedge \clk ) begin
        s492_val_n1 <= s491_val_n1;
    end
    always @(posedge \clk ) begin
        s492_val_n2 <= s491_val_n2;
    end
    always @(posedge \clk ) begin
        s492_val_n3 <= s491_val_n3;
    end
    always @(posedge \clk ) begin
        s492_val_n4 <= s491_val_n4;
    end
    always @(posedge \clk ) begin
        \s493_val  <= \s492_val ;
    end
    always @(posedge \clk ) begin
        s493_val_n1 <= s492_val_n1;
    end
    always @(posedge \clk ) begin
        s493_val_n2 <= s492_val_n2;
    end
    always @(posedge \clk ) begin
        s493_val_n3 <= s492_val_n3;
    end
    always @(posedge \clk ) begin
        s493_val_n4 <= s492_val_n4;
    end
    always @(posedge \clk ) begin
        \s494_val  <= \s493_val ;
    end
    always @(posedge \clk ) begin
        s494_val_n1 <= s493_val_n1;
    end
    always @(posedge \clk ) begin
        s494_val_n2 <= s493_val_n2;
    end
    always @(posedge \clk ) begin
        s494_val_n3 <= s493_val_n3;
    end
    always @(posedge \clk ) begin
        s494_val_n4 <= s493_val_n4;
    end
    always @(posedge \clk ) begin
        \s495_val  <= \s494_val ;
    end
    always @(posedge \clk ) begin
        s495_val_n1 <= s494_val_n1;
    end
    always @(posedge \clk ) begin
        s495_val_n2 <= s494_val_n2;
    end
    always @(posedge \clk ) begin
        s495_val_n3 <= s494_val_n3;
    end
    always @(posedge \clk ) begin
        s495_val_n4 <= s494_val_n4;
    end
    always @(posedge \clk ) begin
        \s496_val  <= \s495_val ;
    end
    always @(posedge \clk ) begin
        s496_val_n1 <= s495_val_n1;
    end
    always @(posedge \clk ) begin
        s496_val_n2 <= s495_val_n2;
    end
    always @(posedge \clk ) begin
        s496_val_n3 <= s495_val_n3;
    end
    always @(posedge \clk ) begin
        s496_val_n4 <= s495_val_n4;
    end
    always @(posedge \clk ) begin
        \s497_val  <= \s496_val ;
    end
    always @(posedge \clk ) begin
        s497_val_n1 <= s496_val_n1;
    end
    always @(posedge \clk ) begin
        s497_val_n2 <= s496_val_n2;
    end
    always @(posedge \clk ) begin
        s497_val_n3 <= s496_val_n3;
    end
    always @(posedge \clk ) begin
        s497_val_n4 <= s496_val_n4;
    end
    always @(posedge \clk ) begin
        \s498_val  <= \s497_val ;
    end
    always @(posedge \clk ) begin
        s498_val_n1 <= s497_val_n1;
    end
    always @(posedge \clk ) begin
        s498_val_n2 <= s497_val_n2;
    end
    always @(posedge \clk ) begin
        s498_val_n3 <= s497_val_n3;
    end
    always @(posedge \clk ) begin
        s498_val_n4 <= s497_val_n4;
    end
    always @(posedge \clk ) begin
        \s499_val  <= \s498_val ;
    end
    always @(posedge \clk ) begin
        s499_val_n1 <= s498_val_n1;
    end
    always @(posedge \clk ) begin
        s499_val_n2 <= s498_val_n2;
    end
    always @(posedge \clk ) begin
        s499_val_n3 <= s498_val_n3;
    end
    always @(posedge \clk ) begin
        s499_val_n4 <= s498_val_n4;
    end
    always @(posedge \clk ) begin
        \s500_val  <= \s499_val ;
    end
    always @(posedge \clk ) begin
        s500_val_n1 <= s499_val_n1;
    end
    always @(posedge \clk ) begin
        s500_val_n2 <= s499_val_n2;
    end
    always @(posedge \clk ) begin
        s500_val_n3 <= s499_val_n3;
    end
    always @(posedge \clk ) begin
        s500_val_n4 <= s499_val_n4;
    end
    always @(posedge \clk ) begin
        \s501_val  <= \s500_val ;
    end
    always @(posedge \clk ) begin
        s501_val_n1 <= s500_val_n1;
    end
    always @(posedge \clk ) begin
        s501_val_n2 <= s500_val_n2;
    end
    always @(posedge \clk ) begin
        s501_val_n3 <= s500_val_n3;
    end
    always @(posedge \clk ) begin
        s501_val_n4 <= s500_val_n4;
    end
    always @(posedge \clk ) begin
        s501_val_n5 <= val_n5;
    end
    always @(posedge \clk ) begin
        \s502_val  <= \s501_val ;
    end
    always @(posedge \clk ) begin
        s502_val_n1 <= s501_val_n1;
    end
    always @(posedge \clk ) begin
        s502_val_n2 <= s501_val_n2;
    end
    always @(posedge \clk ) begin
        s502_val_n3 <= s501_val_n3;
    end
    always @(posedge \clk ) begin
        s502_val_n4 <= s501_val_n4;
    end
    always @(posedge \clk ) begin
        s502_val_n5 <= s501_val_n5;
    end
    always @(posedge \clk ) begin
        \s503_val  <= \s502_val ;
    end
    always @(posedge \clk ) begin
        s503_val_n1 <= s502_val_n1;
    end
    always @(posedge \clk ) begin
        s503_val_n2 <= s502_val_n2;
    end
    always @(posedge \clk ) begin
        s503_val_n3 <= s502_val_n3;
    end
    always @(posedge \clk ) begin
        s503_val_n4 <= s502_val_n4;
    end
    always @(posedge \clk ) begin
        s503_val_n5 <= s502_val_n5;
    end
    always @(posedge \clk ) begin
        \s504_val  <= \s503_val ;
    end
    always @(posedge \clk ) begin
        s504_val_n1 <= s503_val_n1;
    end
    always @(posedge \clk ) begin
        s504_val_n2 <= s503_val_n2;
    end
    always @(posedge \clk ) begin
        s504_val_n3 <= s503_val_n3;
    end
    always @(posedge \clk ) begin
        s504_val_n4 <= s503_val_n4;
    end
    always @(posedge \clk ) begin
        s504_val_n5 <= s503_val_n5;
    end
    always @(posedge \clk ) begin
        \s505_val  <= \s504_val ;
    end
    always @(posedge \clk ) begin
        s505_val_n1 <= s504_val_n1;
    end
    always @(posedge \clk ) begin
        s505_val_n2 <= s504_val_n2;
    end
    always @(posedge \clk ) begin
        s505_val_n3 <= s504_val_n3;
    end
    always @(posedge \clk ) begin
        s505_val_n4 <= s504_val_n4;
    end
    always @(posedge \clk ) begin
        s505_val_n5 <= s504_val_n5;
    end
    always @(posedge \clk ) begin
        \s506_val  <= \s505_val ;
    end
    always @(posedge \clk ) begin
        s506_val_n1 <= s505_val_n1;
    end
    always @(posedge \clk ) begin
        s506_val_n2 <= s505_val_n2;
    end
    always @(posedge \clk ) begin
        s506_val_n3 <= s505_val_n3;
    end
    always @(posedge \clk ) begin
        s506_val_n4 <= s505_val_n4;
    end
    always @(posedge \clk ) begin
        s506_val_n5 <= s505_val_n5;
    end
    always @(posedge \clk ) begin
        \s507_val  <= \s506_val ;
    end
    always @(posedge \clk ) begin
        s507_val_n1 <= s506_val_n1;
    end
    always @(posedge \clk ) begin
        s507_val_n2 <= s506_val_n2;
    end
    always @(posedge \clk ) begin
        s507_val_n3 <= s506_val_n3;
    end
    always @(posedge \clk ) begin
        s507_val_n4 <= s506_val_n4;
    end
    always @(posedge \clk ) begin
        s507_val_n5 <= s506_val_n5;
    end
    always @(posedge \clk ) begin
        \s508_val  <= \s507_val ;
    end
    always @(posedge \clk ) begin
        s508_val_n1 <= s507_val_n1;
    end
    always @(posedge \clk ) begin
        s508_val_n2 <= s507_val_n2;
    end
    always @(posedge \clk ) begin
        s508_val_n3 <= s507_val_n3;
    end
    always @(posedge \clk ) begin
        s508_val_n4 <= s507_val_n4;
    end
    always @(posedge \clk ) begin
        s508_val_n5 <= s507_val_n5;
    end
    always @(posedge \clk ) begin
        \s509_val  <= \s508_val ;
    end
    always @(posedge \clk ) begin
        s509_val_n1 <= s508_val_n1;
    end
    always @(posedge \clk ) begin
        s509_val_n2 <= s508_val_n2;
    end
    always @(posedge \clk ) begin
        s509_val_n3 <= s508_val_n3;
    end
    always @(posedge \clk ) begin
        s509_val_n4 <= s508_val_n4;
    end
    always @(posedge \clk ) begin
        s509_val_n5 <= s508_val_n5;
    end
    always @(posedge \clk ) begin
        \s510_val  <= \s509_val ;
    end
    always @(posedge \clk ) begin
        s510_val_n1 <= s509_val_n1;
    end
    always @(posedge \clk ) begin
        s510_val_n2 <= s509_val_n2;
    end
    always @(posedge \clk ) begin
        s510_val_n3 <= s509_val_n3;
    end
    always @(posedge \clk ) begin
        s510_val_n4 <= s509_val_n4;
    end
    always @(posedge \clk ) begin
        s510_val_n5 <= s509_val_n5;
    end
    always @(posedge \clk ) begin
        \s511_val  <= \s510_val ;
    end
    always @(posedge \clk ) begin
        s511_val_n1 <= s510_val_n1;
    end
    always @(posedge \clk ) begin
        s511_val_n2 <= s510_val_n2;
    end
    always @(posedge \clk ) begin
        s511_val_n3 <= s510_val_n3;
    end
    always @(posedge \clk ) begin
        s511_val_n4 <= s510_val_n4;
    end
    always @(posedge \clk ) begin
        s511_val_n5 <= s510_val_n5;
    end
    always @(posedge \clk ) begin
        \s512_val  <= \s511_val ;
    end
    always @(posedge \clk ) begin
        s512_val_n1 <= s511_val_n1;
    end
    always @(posedge \clk ) begin
        s512_val_n2 <= s511_val_n2;
    end
    always @(posedge \clk ) begin
        s512_val_n3 <= s511_val_n3;
    end
    always @(posedge \clk ) begin
        s512_val_n4 <= s511_val_n4;
    end
    always @(posedge \clk ) begin
        s512_val_n5 <= s511_val_n5;
    end
    always @(posedge \clk ) begin
        \s513_val  <= \s512_val ;
    end
    always @(posedge \clk ) begin
        s513_val_n1 <= s512_val_n1;
    end
    always @(posedge \clk ) begin
        s513_val_n2 <= s512_val_n2;
    end
    always @(posedge \clk ) begin
        s513_val_n3 <= s512_val_n3;
    end
    always @(posedge \clk ) begin
        s513_val_n4 <= s512_val_n4;
    end
    always @(posedge \clk ) begin
        s513_val_n5 <= s512_val_n5;
    end
    always @(posedge \clk ) begin
        \s514_val  <= \s513_val ;
    end
    always @(posedge \clk ) begin
        s514_val_n1 <= s513_val_n1;
    end
    always @(posedge \clk ) begin
        s514_val_n2 <= s513_val_n2;
    end
    always @(posedge \clk ) begin
        s514_val_n3 <= s513_val_n3;
    end
    always @(posedge \clk ) begin
        s514_val_n4 <= s513_val_n4;
    end
    always @(posedge \clk ) begin
        s514_val_n5 <= s513_val_n5;
    end
    always @(posedge \clk ) begin
        \s515_val  <= \s514_val ;
    end
    always @(posedge \clk ) begin
        s515_val_n1 <= s514_val_n1;
    end
    always @(posedge \clk ) begin
        s515_val_n2 <= s514_val_n2;
    end
    always @(posedge \clk ) begin
        s515_val_n3 <= s514_val_n3;
    end
    always @(posedge \clk ) begin
        s515_val_n4 <= s514_val_n4;
    end
    always @(posedge \clk ) begin
        s515_val_n5 <= s514_val_n5;
    end
    always @(posedge \clk ) begin
        \s516_val  <= \s515_val ;
    end
    always @(posedge \clk ) begin
        s516_val_n1 <= s515_val_n1;
    end
    always @(posedge \clk ) begin
        s516_val_n2 <= s515_val_n2;
    end
    always @(posedge \clk ) begin
        s516_val_n3 <= s515_val_n3;
    end
    always @(posedge \clk ) begin
        s516_val_n4 <= s515_val_n4;
    end
    always @(posedge \clk ) begin
        s516_val_n5 <= s515_val_n5;
    end
    always @(posedge \clk ) begin
        \s517_val  <= \s516_val ;
    end
    always @(posedge \clk ) begin
        s517_val_n1 <= s516_val_n1;
    end
    always @(posedge \clk ) begin
        s517_val_n2 <= s516_val_n2;
    end
    always @(posedge \clk ) begin
        s517_val_n3 <= s516_val_n3;
    end
    always @(posedge \clk ) begin
        s517_val_n4 <= s516_val_n4;
    end
    always @(posedge \clk ) begin
        s517_val_n5 <= s516_val_n5;
    end
    always @(posedge \clk ) begin
        \s518_val  <= \s517_val ;
    end
    always @(posedge \clk ) begin
        s518_val_n1 <= s517_val_n1;
    end
    always @(posedge \clk ) begin
        s518_val_n2 <= s517_val_n2;
    end
    always @(posedge \clk ) begin
        s518_val_n3 <= s517_val_n3;
    end
    always @(posedge \clk ) begin
        s518_val_n4 <= s517_val_n4;
    end
    always @(posedge \clk ) begin
        s518_val_n5 <= s517_val_n5;
    end
    always @(posedge \clk ) begin
        \s519_val  <= \s518_val ;
    end
    always @(posedge \clk ) begin
        s519_val_n1 <= s518_val_n1;
    end
    always @(posedge \clk ) begin
        s519_val_n2 <= s518_val_n2;
    end
    always @(posedge \clk ) begin
        s519_val_n3 <= s518_val_n3;
    end
    always @(posedge \clk ) begin
        s519_val_n4 <= s518_val_n4;
    end
    always @(posedge \clk ) begin
        s519_val_n5 <= s518_val_n5;
    end
    always @(posedge \clk ) begin
        \s520_val  <= \s519_val ;
    end
    always @(posedge \clk ) begin
        s520_val_n1 <= s519_val_n1;
    end
    always @(posedge \clk ) begin
        s520_val_n2 <= s519_val_n2;
    end
    always @(posedge \clk ) begin
        s520_val_n3 <= s519_val_n3;
    end
    always @(posedge \clk ) begin
        s520_val_n4 <= s519_val_n4;
    end
    always @(posedge \clk ) begin
        s520_val_n5 <= s519_val_n5;
    end
    always @(posedge \clk ) begin
        \s521_val  <= \s520_val ;
    end
    always @(posedge \clk ) begin
        s521_val_n1 <= s520_val_n1;
    end
    always @(posedge \clk ) begin
        s521_val_n2 <= s520_val_n2;
    end
    always @(posedge \clk ) begin
        s521_val_n3 <= s520_val_n3;
    end
    always @(posedge \clk ) begin
        s521_val_n4 <= s520_val_n4;
    end
    always @(posedge \clk ) begin
        s521_val_n5 <= s520_val_n5;
    end
    always @(posedge \clk ) begin
        \s522_val  <= \s521_val ;
    end
    always @(posedge \clk ) begin
        s522_val_n1 <= s521_val_n1;
    end
    always @(posedge \clk ) begin
        s522_val_n2 <= s521_val_n2;
    end
    always @(posedge \clk ) begin
        s522_val_n3 <= s521_val_n3;
    end
    always @(posedge \clk ) begin
        s522_val_n4 <= s521_val_n4;
    end
    always @(posedge \clk ) begin
        s522_val_n5 <= s521_val_n5;
    end
    always @(posedge \clk ) begin
        \s523_val  <= \s522_val ;
    end
    always @(posedge \clk ) begin
        s523_val_n1 <= s522_val_n1;
    end
    always @(posedge \clk ) begin
        s523_val_n2 <= s522_val_n2;
    end
    always @(posedge \clk ) begin
        s523_val_n3 <= s522_val_n3;
    end
    always @(posedge \clk ) begin
        s523_val_n4 <= s522_val_n4;
    end
    always @(posedge \clk ) begin
        s523_val_n5 <= s522_val_n5;
    end
    always @(posedge \clk ) begin
        \s524_val  <= \s523_val ;
    end
    always @(posedge \clk ) begin
        s524_val_n1 <= s523_val_n1;
    end
    always @(posedge \clk ) begin
        s524_val_n2 <= s523_val_n2;
    end
    always @(posedge \clk ) begin
        s524_val_n3 <= s523_val_n3;
    end
    always @(posedge \clk ) begin
        s524_val_n4 <= s523_val_n4;
    end
    always @(posedge \clk ) begin
        s524_val_n5 <= s523_val_n5;
    end
    always @(posedge \clk ) begin
        \s525_val  <= \s524_val ;
    end
    always @(posedge \clk ) begin
        s525_val_n1 <= s524_val_n1;
    end
    always @(posedge \clk ) begin
        s525_val_n2 <= s524_val_n2;
    end
    always @(posedge \clk ) begin
        s525_val_n3 <= s524_val_n3;
    end
    always @(posedge \clk ) begin
        s525_val_n4 <= s524_val_n4;
    end
    always @(posedge \clk ) begin
        s525_val_n5 <= s524_val_n5;
    end
    always @(posedge \clk ) begin
        \s526_val  <= \s525_val ;
    end
    always @(posedge \clk ) begin
        s526_val_n1 <= s525_val_n1;
    end
    always @(posedge \clk ) begin
        s526_val_n2 <= s525_val_n2;
    end
    always @(posedge \clk ) begin
        s526_val_n3 <= s525_val_n3;
    end
    always @(posedge \clk ) begin
        s526_val_n4 <= s525_val_n4;
    end
    always @(posedge \clk ) begin
        s526_val_n5 <= s525_val_n5;
    end
    always @(posedge \clk ) begin
        \s527_val  <= \s526_val ;
    end
    always @(posedge \clk ) begin
        s527_val_n1 <= s526_val_n1;
    end
    always @(posedge \clk ) begin
        s527_val_n2 <= s526_val_n2;
    end
    always @(posedge \clk ) begin
        s527_val_n3 <= s526_val_n3;
    end
    always @(posedge \clk ) begin
        s527_val_n4 <= s526_val_n4;
    end
    always @(posedge \clk ) begin
        s527_val_n5 <= s526_val_n5;
    end
    always @(posedge \clk ) begin
        \s528_val  <= \s527_val ;
    end
    always @(posedge \clk ) begin
        s528_val_n1 <= s527_val_n1;
    end
    always @(posedge \clk ) begin
        s528_val_n2 <= s527_val_n2;
    end
    always @(posedge \clk ) begin
        s528_val_n3 <= s527_val_n3;
    end
    always @(posedge \clk ) begin
        s528_val_n4 <= s527_val_n4;
    end
    always @(posedge \clk ) begin
        s528_val_n5 <= s527_val_n5;
    end
    always @(posedge \clk ) begin
        \s529_val  <= \s528_val ;
    end
    always @(posedge \clk ) begin
        s529_val_n1 <= s528_val_n1;
    end
    always @(posedge \clk ) begin
        s529_val_n2 <= s528_val_n2;
    end
    always @(posedge \clk ) begin
        s529_val_n3 <= s528_val_n3;
    end
    always @(posedge \clk ) begin
        s529_val_n4 <= s528_val_n4;
    end
    always @(posedge \clk ) begin
        s529_val_n5 <= s528_val_n5;
    end
    always @(posedge \clk ) begin
        \s530_val  <= \s529_val ;
    end
    always @(posedge \clk ) begin
        s530_val_n1 <= s529_val_n1;
    end
    always @(posedge \clk ) begin
        s530_val_n2 <= s529_val_n2;
    end
    always @(posedge \clk ) begin
        s530_val_n3 <= s529_val_n3;
    end
    always @(posedge \clk ) begin
        s530_val_n4 <= s529_val_n4;
    end
    always @(posedge \clk ) begin
        s530_val_n5 <= s529_val_n5;
    end
    always @(posedge \clk ) begin
        \s531_val  <= \s530_val ;
    end
    always @(posedge \clk ) begin
        s531_val_n1 <= s530_val_n1;
    end
    always @(posedge \clk ) begin
        s531_val_n2 <= s530_val_n2;
    end
    always @(posedge \clk ) begin
        s531_val_n3 <= s530_val_n3;
    end
    always @(posedge \clk ) begin
        s531_val_n4 <= s530_val_n4;
    end
    always @(posedge \clk ) begin
        s531_val_n5 <= s530_val_n5;
    end
    always @(posedge \clk ) begin
        \s532_val  <= \s531_val ;
    end
    always @(posedge \clk ) begin
        s532_val_n1 <= s531_val_n1;
    end
    always @(posedge \clk ) begin
        s532_val_n2 <= s531_val_n2;
    end
    always @(posedge \clk ) begin
        s532_val_n3 <= s531_val_n3;
    end
    always @(posedge \clk ) begin
        s532_val_n4 <= s531_val_n4;
    end
    always @(posedge \clk ) begin
        s532_val_n5 <= s531_val_n5;
    end
    always @(posedge \clk ) begin
        \s533_val  <= \s532_val ;
    end
    always @(posedge \clk ) begin
        s533_val_n1 <= s532_val_n1;
    end
    always @(posedge \clk ) begin
        s533_val_n2 <= s532_val_n2;
    end
    always @(posedge \clk ) begin
        s533_val_n3 <= s532_val_n3;
    end
    always @(posedge \clk ) begin
        s533_val_n4 <= s532_val_n4;
    end
    always @(posedge \clk ) begin
        s533_val_n5 <= s532_val_n5;
    end
    always @(posedge \clk ) begin
        \s534_val  <= \s533_val ;
    end
    always @(posedge \clk ) begin
        s534_val_n1 <= s533_val_n1;
    end
    always @(posedge \clk ) begin
        s534_val_n2 <= s533_val_n2;
    end
    always @(posedge \clk ) begin
        s534_val_n3 <= s533_val_n3;
    end
    always @(posedge \clk ) begin
        s534_val_n4 <= s533_val_n4;
    end
    always @(posedge \clk ) begin
        s534_val_n5 <= s533_val_n5;
    end
    always @(posedge \clk ) begin
        \s535_val  <= \s534_val ;
    end
    always @(posedge \clk ) begin
        s535_val_n1 <= s534_val_n1;
    end
    always @(posedge \clk ) begin
        s535_val_n2 <= s534_val_n2;
    end
    always @(posedge \clk ) begin
        s535_val_n3 <= s534_val_n3;
    end
    always @(posedge \clk ) begin
        s535_val_n4 <= s534_val_n4;
    end
    always @(posedge \clk ) begin
        s535_val_n5 <= s534_val_n5;
    end
    always @(posedge \clk ) begin
        \s536_val  <= \s535_val ;
    end
    always @(posedge \clk ) begin
        s536_val_n1 <= s535_val_n1;
    end
    always @(posedge \clk ) begin
        s536_val_n2 <= s535_val_n2;
    end
    always @(posedge \clk ) begin
        s536_val_n3 <= s535_val_n3;
    end
    always @(posedge \clk ) begin
        s536_val_n4 <= s535_val_n4;
    end
    always @(posedge \clk ) begin
        s536_val_n5 <= s535_val_n5;
    end
    always @(posedge \clk ) begin
        \s537_val  <= \s536_val ;
    end
    always @(posedge \clk ) begin
        s537_val_n1 <= s536_val_n1;
    end
    always @(posedge \clk ) begin
        s537_val_n2 <= s536_val_n2;
    end
    always @(posedge \clk ) begin
        s537_val_n3 <= s536_val_n3;
    end
    always @(posedge \clk ) begin
        s537_val_n4 <= s536_val_n4;
    end
    always @(posedge \clk ) begin
        s537_val_n5 <= s536_val_n5;
    end
    always @(posedge \clk ) begin
        \s538_val  <= \s537_val ;
    end
    always @(posedge \clk ) begin
        s538_val_n1 <= s537_val_n1;
    end
    always @(posedge \clk ) begin
        s538_val_n2 <= s537_val_n2;
    end
    always @(posedge \clk ) begin
        s538_val_n3 <= s537_val_n3;
    end
    always @(posedge \clk ) begin
        s538_val_n4 <= s537_val_n4;
    end
    always @(posedge \clk ) begin
        s538_val_n5 <= s537_val_n5;
    end
    always @(posedge \clk ) begin
        \s539_val  <= \s538_val ;
    end
    always @(posedge \clk ) begin
        s539_val_n1 <= s538_val_n1;
    end
    always @(posedge \clk ) begin
        s539_val_n2 <= s538_val_n2;
    end
    always @(posedge \clk ) begin
        s539_val_n3 <= s538_val_n3;
    end
    always @(posedge \clk ) begin
        s539_val_n4 <= s538_val_n4;
    end
    always @(posedge \clk ) begin
        s539_val_n5 <= s538_val_n5;
    end
    always @(posedge \clk ) begin
        \s540_val  <= \s539_val ;
    end
    always @(posedge \clk ) begin
        s540_val_n1 <= s539_val_n1;
    end
    always @(posedge \clk ) begin
        s540_val_n2 <= s539_val_n2;
    end
    always @(posedge \clk ) begin
        s540_val_n3 <= s539_val_n3;
    end
    always @(posedge \clk ) begin
        s540_val_n4 <= s539_val_n4;
    end
    always @(posedge \clk ) begin
        s540_val_n5 <= s539_val_n5;
    end
    always @(posedge \clk ) begin
        \s541_val  <= \s540_val ;
    end
    always @(posedge \clk ) begin
        s541_val_n1 <= s540_val_n1;
    end
    always @(posedge \clk ) begin
        s541_val_n2 <= s540_val_n2;
    end
    always @(posedge \clk ) begin
        s541_val_n3 <= s540_val_n3;
    end
    always @(posedge \clk ) begin
        s541_val_n4 <= s540_val_n4;
    end
    always @(posedge \clk ) begin
        s541_val_n5 <= s540_val_n5;
    end
    always @(posedge \clk ) begin
        \s542_val  <= \s541_val ;
    end
    always @(posedge \clk ) begin
        s542_val_n1 <= s541_val_n1;
    end
    always @(posedge \clk ) begin
        s542_val_n2 <= s541_val_n2;
    end
    always @(posedge \clk ) begin
        s542_val_n3 <= s541_val_n3;
    end
    always @(posedge \clk ) begin
        s542_val_n4 <= s541_val_n4;
    end
    always @(posedge \clk ) begin
        s542_val_n5 <= s541_val_n5;
    end
    always @(posedge \clk ) begin
        \s543_val  <= \s542_val ;
    end
    always @(posedge \clk ) begin
        s543_val_n1 <= s542_val_n1;
    end
    always @(posedge \clk ) begin
        s543_val_n2 <= s542_val_n2;
    end
    always @(posedge \clk ) begin
        s543_val_n3 <= s542_val_n3;
    end
    always @(posedge \clk ) begin
        s543_val_n4 <= s542_val_n4;
    end
    always @(posedge \clk ) begin
        s543_val_n5 <= s542_val_n5;
    end
    always @(posedge \clk ) begin
        \s544_val  <= \s543_val ;
    end
    always @(posedge \clk ) begin
        s544_val_n1 <= s543_val_n1;
    end
    always @(posedge \clk ) begin
        s544_val_n2 <= s543_val_n2;
    end
    always @(posedge \clk ) begin
        s544_val_n3 <= s543_val_n3;
    end
    always @(posedge \clk ) begin
        s544_val_n4 <= s543_val_n4;
    end
    always @(posedge \clk ) begin
        s544_val_n5 <= s543_val_n5;
    end
    always @(posedge \clk ) begin
        \s545_val  <= \s544_val ;
    end
    always @(posedge \clk ) begin
        s545_val_n1 <= s544_val_n1;
    end
    always @(posedge \clk ) begin
        s545_val_n2 <= s544_val_n2;
    end
    always @(posedge \clk ) begin
        s545_val_n3 <= s544_val_n3;
    end
    always @(posedge \clk ) begin
        s545_val_n4 <= s544_val_n4;
    end
    always @(posedge \clk ) begin
        s545_val_n5 <= s544_val_n5;
    end
    always @(posedge \clk ) begin
        \s546_val  <= \s545_val ;
    end
    always @(posedge \clk ) begin
        s546_val_n1 <= s545_val_n1;
    end
    always @(posedge \clk ) begin
        s546_val_n2 <= s545_val_n2;
    end
    always @(posedge \clk ) begin
        s546_val_n3 <= s545_val_n3;
    end
    always @(posedge \clk ) begin
        s546_val_n4 <= s545_val_n4;
    end
    always @(posedge \clk ) begin
        s546_val_n5 <= s545_val_n5;
    end
    always @(posedge \clk ) begin
        \s547_val  <= \s546_val ;
    end
    always @(posedge \clk ) begin
        s547_val_n1 <= s546_val_n1;
    end
    always @(posedge \clk ) begin
        s547_val_n2 <= s546_val_n2;
    end
    always @(posedge \clk ) begin
        s547_val_n3 <= s546_val_n3;
    end
    always @(posedge \clk ) begin
        s547_val_n4 <= s546_val_n4;
    end
    always @(posedge \clk ) begin
        s547_val_n5 <= s546_val_n5;
    end
    always @(posedge \clk ) begin
        \s548_val  <= \s547_val ;
    end
    always @(posedge \clk ) begin
        s548_val_n1 <= s547_val_n1;
    end
    always @(posedge \clk ) begin
        s548_val_n2 <= s547_val_n2;
    end
    always @(posedge \clk ) begin
        s548_val_n3 <= s547_val_n3;
    end
    always @(posedge \clk ) begin
        s548_val_n4 <= s547_val_n4;
    end
    always @(posedge \clk ) begin
        s548_val_n5 <= s547_val_n5;
    end
    always @(posedge \clk ) begin
        \s549_val  <= \s548_val ;
    end
    always @(posedge \clk ) begin
        s549_val_n1 <= s548_val_n1;
    end
    always @(posedge \clk ) begin
        s549_val_n2 <= s548_val_n2;
    end
    always @(posedge \clk ) begin
        s549_val_n3 <= s548_val_n3;
    end
    always @(posedge \clk ) begin
        s549_val_n4 <= s548_val_n4;
    end
    always @(posedge \clk ) begin
        s549_val_n5 <= s548_val_n5;
    end
    always @(posedge \clk ) begin
        \s550_val  <= \s549_val ;
    end
    always @(posedge \clk ) begin
        s550_val_n1 <= s549_val_n1;
    end
    always @(posedge \clk ) begin
        s550_val_n2 <= s549_val_n2;
    end
    always @(posedge \clk ) begin
        s550_val_n3 <= s549_val_n3;
    end
    always @(posedge \clk ) begin
        s550_val_n4 <= s549_val_n4;
    end
    always @(posedge \clk ) begin
        s550_val_n5 <= s549_val_n5;
    end
    always @(posedge \clk ) begin
        \s551_val  <= \s550_val ;
    end
    always @(posedge \clk ) begin
        s551_val_n1 <= s550_val_n1;
    end
    always @(posedge \clk ) begin
        s551_val_n2 <= s550_val_n2;
    end
    always @(posedge \clk ) begin
        s551_val_n3 <= s550_val_n3;
    end
    always @(posedge \clk ) begin
        s551_val_n4 <= s550_val_n4;
    end
    always @(posedge \clk ) begin
        s551_val_n5 <= s550_val_n5;
    end
    always @(posedge \clk ) begin
        \s552_val  <= \s551_val ;
    end
    always @(posedge \clk ) begin
        s552_val_n1 <= s551_val_n1;
    end
    always @(posedge \clk ) begin
        s552_val_n2 <= s551_val_n2;
    end
    always @(posedge \clk ) begin
        s552_val_n3 <= s551_val_n3;
    end
    always @(posedge \clk ) begin
        s552_val_n4 <= s551_val_n4;
    end
    always @(posedge \clk ) begin
        s552_val_n5 <= s551_val_n5;
    end
    always @(posedge \clk ) begin
        \s553_val  <= \s552_val ;
    end
    always @(posedge \clk ) begin
        s553_val_n1 <= s552_val_n1;
    end
    always @(posedge \clk ) begin
        s553_val_n2 <= s552_val_n2;
    end
    always @(posedge \clk ) begin
        s553_val_n3 <= s552_val_n3;
    end
    always @(posedge \clk ) begin
        s553_val_n4 <= s552_val_n4;
    end
    always @(posedge \clk ) begin
        s553_val_n5 <= s552_val_n5;
    end
    always @(posedge \clk ) begin
        \s554_val  <= \s553_val ;
    end
    always @(posedge \clk ) begin
        s554_val_n1 <= s553_val_n1;
    end
    always @(posedge \clk ) begin
        s554_val_n2 <= s553_val_n2;
    end
    always @(posedge \clk ) begin
        s554_val_n3 <= s553_val_n3;
    end
    always @(posedge \clk ) begin
        s554_val_n4 <= s553_val_n4;
    end
    always @(posedge \clk ) begin
        s554_val_n5 <= s553_val_n5;
    end
    always @(posedge \clk ) begin
        \s555_val  <= \s554_val ;
    end
    always @(posedge \clk ) begin
        s555_val_n1 <= s554_val_n1;
    end
    always @(posedge \clk ) begin
        s555_val_n2 <= s554_val_n2;
    end
    always @(posedge \clk ) begin
        s555_val_n3 <= s554_val_n3;
    end
    always @(posedge \clk ) begin
        s555_val_n4 <= s554_val_n4;
    end
    always @(posedge \clk ) begin
        s555_val_n5 <= s554_val_n5;
    end
    always @(posedge \clk ) begin
        \s556_val  <= \s555_val ;
    end
    always @(posedge \clk ) begin
        s556_val_n1 <= s555_val_n1;
    end
    always @(posedge \clk ) begin
        s556_val_n2 <= s555_val_n2;
    end
    always @(posedge \clk ) begin
        s556_val_n3 <= s555_val_n3;
    end
    always @(posedge \clk ) begin
        s556_val_n4 <= s555_val_n4;
    end
    always @(posedge \clk ) begin
        s556_val_n5 <= s555_val_n5;
    end
    always @(posedge \clk ) begin
        \s557_val  <= \s556_val ;
    end
    always @(posedge \clk ) begin
        s557_val_n1 <= s556_val_n1;
    end
    always @(posedge \clk ) begin
        s557_val_n2 <= s556_val_n2;
    end
    always @(posedge \clk ) begin
        s557_val_n3 <= s556_val_n3;
    end
    always @(posedge \clk ) begin
        s557_val_n4 <= s556_val_n4;
    end
    always @(posedge \clk ) begin
        s557_val_n5 <= s556_val_n5;
    end
    always @(posedge \clk ) begin
        \s558_val  <= \s557_val ;
    end
    always @(posedge \clk ) begin
        s558_val_n1 <= s557_val_n1;
    end
    always @(posedge \clk ) begin
        s558_val_n2 <= s557_val_n2;
    end
    always @(posedge \clk ) begin
        s558_val_n3 <= s557_val_n3;
    end
    always @(posedge \clk ) begin
        s558_val_n4 <= s557_val_n4;
    end
    always @(posedge \clk ) begin
        s558_val_n5 <= s557_val_n5;
    end
    always @(posedge \clk ) begin
        \s559_val  <= \s558_val ;
    end
    always @(posedge \clk ) begin
        s559_val_n1 <= s558_val_n1;
    end
    always @(posedge \clk ) begin
        s559_val_n2 <= s558_val_n2;
    end
    always @(posedge \clk ) begin
        s559_val_n3 <= s558_val_n3;
    end
    always @(posedge \clk ) begin
        s559_val_n4 <= s558_val_n4;
    end
    always @(posedge \clk ) begin
        s559_val_n5 <= s558_val_n5;
    end
    always @(posedge \clk ) begin
        \s560_val  <= \s559_val ;
    end
    always @(posedge \clk ) begin
        s560_val_n1 <= s559_val_n1;
    end
    always @(posedge \clk ) begin
        s560_val_n2 <= s559_val_n2;
    end
    always @(posedge \clk ) begin
        s560_val_n3 <= s559_val_n3;
    end
    always @(posedge \clk ) begin
        s560_val_n4 <= s559_val_n4;
    end
    always @(posedge \clk ) begin
        s560_val_n5 <= s559_val_n5;
    end
    always @(posedge \clk ) begin
        \s561_val  <= \s560_val ;
    end
    always @(posedge \clk ) begin
        s561_val_n1 <= s560_val_n1;
    end
    always @(posedge \clk ) begin
        s561_val_n2 <= s560_val_n2;
    end
    always @(posedge \clk ) begin
        s561_val_n3 <= s560_val_n3;
    end
    always @(posedge \clk ) begin
        s561_val_n4 <= s560_val_n4;
    end
    always @(posedge \clk ) begin
        s561_val_n5 <= s560_val_n5;
    end
    always @(posedge \clk ) begin
        \s562_val  <= \s561_val ;
    end
    always @(posedge \clk ) begin
        s562_val_n1 <= s561_val_n1;
    end
    always @(posedge \clk ) begin
        s562_val_n2 <= s561_val_n2;
    end
    always @(posedge \clk ) begin
        s562_val_n3 <= s561_val_n3;
    end
    always @(posedge \clk ) begin
        s562_val_n4 <= s561_val_n4;
    end
    always @(posedge \clk ) begin
        s562_val_n5 <= s561_val_n5;
    end
    always @(posedge \clk ) begin
        \s563_val  <= \s562_val ;
    end
    always @(posedge \clk ) begin
        s563_val_n1 <= s562_val_n1;
    end
    always @(posedge \clk ) begin
        s563_val_n2 <= s562_val_n2;
    end
    always @(posedge \clk ) begin
        s563_val_n3 <= s562_val_n3;
    end
    always @(posedge \clk ) begin
        s563_val_n4 <= s562_val_n4;
    end
    always @(posedge \clk ) begin
        s563_val_n5 <= s562_val_n5;
    end
    always @(posedge \clk ) begin
        \s564_val  <= \s563_val ;
    end
    always @(posedge \clk ) begin
        s564_val_n1 <= s563_val_n1;
    end
    always @(posedge \clk ) begin
        s564_val_n2 <= s563_val_n2;
    end
    always @(posedge \clk ) begin
        s564_val_n3 <= s563_val_n3;
    end
    always @(posedge \clk ) begin
        s564_val_n4 <= s563_val_n4;
    end
    always @(posedge \clk ) begin
        s564_val_n5 <= s563_val_n5;
    end
    always @(posedge \clk ) begin
        \s565_val  <= \s564_val ;
    end
    always @(posedge \clk ) begin
        s565_val_n1 <= s564_val_n1;
    end
    always @(posedge \clk ) begin
        s565_val_n2 <= s564_val_n2;
    end
    always @(posedge \clk ) begin
        s565_val_n3 <= s564_val_n3;
    end
    always @(posedge \clk ) begin
        s565_val_n4 <= s564_val_n4;
    end
    always @(posedge \clk ) begin
        s565_val_n5 <= s564_val_n5;
    end
    always @(posedge \clk ) begin
        \s566_val  <= \s565_val ;
    end
    always @(posedge \clk ) begin
        s566_val_n1 <= s565_val_n1;
    end
    always @(posedge \clk ) begin
        s566_val_n2 <= s565_val_n2;
    end
    always @(posedge \clk ) begin
        s566_val_n3 <= s565_val_n3;
    end
    always @(posedge \clk ) begin
        s566_val_n4 <= s565_val_n4;
    end
    always @(posedge \clk ) begin
        s566_val_n5 <= s565_val_n5;
    end
    always @(posedge \clk ) begin
        \s567_val  <= \s566_val ;
    end
    always @(posedge \clk ) begin
        s567_val_n1 <= s566_val_n1;
    end
    always @(posedge \clk ) begin
        s567_val_n2 <= s566_val_n2;
    end
    always @(posedge \clk ) begin
        s567_val_n3 <= s566_val_n3;
    end
    always @(posedge \clk ) begin
        s567_val_n4 <= s566_val_n4;
    end
    always @(posedge \clk ) begin
        s567_val_n5 <= s566_val_n5;
    end
    always @(posedge \clk ) begin
        \s568_val  <= \s567_val ;
    end
    always @(posedge \clk ) begin
        s568_val_n1 <= s567_val_n1;
    end
    always @(posedge \clk ) begin
        s568_val_n2 <= s567_val_n2;
    end
    always @(posedge \clk ) begin
        s568_val_n3 <= s567_val_n3;
    end
    always @(posedge \clk ) begin
        s568_val_n4 <= s567_val_n4;
    end
    always @(posedge \clk ) begin
        s568_val_n5 <= s567_val_n5;
    end
    always @(posedge \clk ) begin
        \s569_val  <= \s568_val ;
    end
    always @(posedge \clk ) begin
        s569_val_n1 <= s568_val_n1;
    end
    always @(posedge \clk ) begin
        s569_val_n2 <= s568_val_n2;
    end
    always @(posedge \clk ) begin
        s569_val_n3 <= s568_val_n3;
    end
    always @(posedge \clk ) begin
        s569_val_n4 <= s568_val_n4;
    end
    always @(posedge \clk ) begin
        s569_val_n5 <= s568_val_n5;
    end
    always @(posedge \clk ) begin
        \s570_val  <= \s569_val ;
    end
    always @(posedge \clk ) begin
        s570_val_n1 <= s569_val_n1;
    end
    always @(posedge \clk ) begin
        s570_val_n2 <= s569_val_n2;
    end
    always @(posedge \clk ) begin
        s570_val_n3 <= s569_val_n3;
    end
    always @(posedge \clk ) begin
        s570_val_n4 <= s569_val_n4;
    end
    always @(posedge \clk ) begin
        s570_val_n5 <= s569_val_n5;
    end
    always @(posedge \clk ) begin
        \s571_val  <= \s570_val ;
    end
    always @(posedge \clk ) begin
        s571_val_n1 <= s570_val_n1;
    end
    always @(posedge \clk ) begin
        s571_val_n2 <= s570_val_n2;
    end
    always @(posedge \clk ) begin
        s571_val_n3 <= s570_val_n3;
    end
    always @(posedge \clk ) begin
        s571_val_n4 <= s570_val_n4;
    end
    always @(posedge \clk ) begin
        s571_val_n5 <= s570_val_n5;
    end
    always @(posedge \clk ) begin
        \s572_val  <= \s571_val ;
    end
    always @(posedge \clk ) begin
        s572_val_n1 <= s571_val_n1;
    end
    always @(posedge \clk ) begin
        s572_val_n2 <= s571_val_n2;
    end
    always @(posedge \clk ) begin
        s572_val_n3 <= s571_val_n3;
    end
    always @(posedge \clk ) begin
        s572_val_n4 <= s571_val_n4;
    end
    always @(posedge \clk ) begin
        s572_val_n5 <= s571_val_n5;
    end
    always @(posedge \clk ) begin
        \s573_val  <= \s572_val ;
    end
    always @(posedge \clk ) begin
        s573_val_n1 <= s572_val_n1;
    end
    always @(posedge \clk ) begin
        s573_val_n2 <= s572_val_n2;
    end
    always @(posedge \clk ) begin
        s573_val_n3 <= s572_val_n3;
    end
    always @(posedge \clk ) begin
        s573_val_n4 <= s572_val_n4;
    end
    always @(posedge \clk ) begin
        s573_val_n5 <= s572_val_n5;
    end
    always @(posedge \clk ) begin
        \s574_val  <= \s573_val ;
    end
    always @(posedge \clk ) begin
        s574_val_n1 <= s573_val_n1;
    end
    always @(posedge \clk ) begin
        s574_val_n2 <= s573_val_n2;
    end
    always @(posedge \clk ) begin
        s574_val_n3 <= s573_val_n3;
    end
    always @(posedge \clk ) begin
        s574_val_n4 <= s573_val_n4;
    end
    always @(posedge \clk ) begin
        s574_val_n5 <= s573_val_n5;
    end
    always @(posedge \clk ) begin
        \s575_val  <= \s574_val ;
    end
    always @(posedge \clk ) begin
        s575_val_n1 <= s574_val_n1;
    end
    always @(posedge \clk ) begin
        s575_val_n2 <= s574_val_n2;
    end
    always @(posedge \clk ) begin
        s575_val_n3 <= s574_val_n3;
    end
    always @(posedge \clk ) begin
        s575_val_n4 <= s574_val_n4;
    end
    always @(posedge \clk ) begin
        s575_val_n5 <= s574_val_n5;
    end
    always @(posedge \clk ) begin
        \s576_val  <= \s575_val ;
    end
    always @(posedge \clk ) begin
        s576_val_n1 <= s575_val_n1;
    end
    always @(posedge \clk ) begin
        s576_val_n2 <= s575_val_n2;
    end
    always @(posedge \clk ) begin
        s576_val_n3 <= s575_val_n3;
    end
    always @(posedge \clk ) begin
        s576_val_n4 <= s575_val_n4;
    end
    always @(posedge \clk ) begin
        s576_val_n5 <= s575_val_n5;
    end
    always @(posedge \clk ) begin
        \s577_val  <= \s576_val ;
    end
    always @(posedge \clk ) begin
        s577_val_n1 <= s576_val_n1;
    end
    always @(posedge \clk ) begin
        s577_val_n2 <= s576_val_n2;
    end
    always @(posedge \clk ) begin
        s577_val_n3 <= s576_val_n3;
    end
    always @(posedge \clk ) begin
        s577_val_n4 <= s576_val_n4;
    end
    always @(posedge \clk ) begin
        s577_val_n5 <= s576_val_n5;
    end
    always @(posedge \clk ) begin
        \s578_val  <= \s577_val ;
    end
    always @(posedge \clk ) begin
        s578_val_n1 <= s577_val_n1;
    end
    always @(posedge \clk ) begin
        s578_val_n2 <= s577_val_n2;
    end
    always @(posedge \clk ) begin
        s578_val_n3 <= s577_val_n3;
    end
    always @(posedge \clk ) begin
        s578_val_n4 <= s577_val_n4;
    end
    always @(posedge \clk ) begin
        s578_val_n5 <= s577_val_n5;
    end
    always @(posedge \clk ) begin
        \s579_val  <= \s578_val ;
    end
    always @(posedge \clk ) begin
        s579_val_n1 <= s578_val_n1;
    end
    always @(posedge \clk ) begin
        s579_val_n2 <= s578_val_n2;
    end
    always @(posedge \clk ) begin
        s579_val_n3 <= s578_val_n3;
    end
    always @(posedge \clk ) begin
        s579_val_n4 <= s578_val_n4;
    end
    always @(posedge \clk ) begin
        s579_val_n5 <= s578_val_n5;
    end
    always @(posedge \clk ) begin
        \s580_val  <= \s579_val ;
    end
    always @(posedge \clk ) begin
        s580_val_n1 <= s579_val_n1;
    end
    always @(posedge \clk ) begin
        s580_val_n2 <= s579_val_n2;
    end
    always @(posedge \clk ) begin
        s580_val_n3 <= s579_val_n3;
    end
    always @(posedge \clk ) begin
        s580_val_n4 <= s579_val_n4;
    end
    always @(posedge \clk ) begin
        s580_val_n5 <= s579_val_n5;
    end
    always @(posedge \clk ) begin
        \s581_val  <= \s580_val ;
    end
    always @(posedge \clk ) begin
        s581_val_n1 <= s580_val_n1;
    end
    always @(posedge \clk ) begin
        s581_val_n2 <= s580_val_n2;
    end
    always @(posedge \clk ) begin
        s581_val_n3 <= s580_val_n3;
    end
    always @(posedge \clk ) begin
        s581_val_n4 <= s580_val_n4;
    end
    always @(posedge \clk ) begin
        s581_val_n5 <= s580_val_n5;
    end
    always @(posedge \clk ) begin
        \s582_val  <= \s581_val ;
    end
    always @(posedge \clk ) begin
        s582_val_n1 <= s581_val_n1;
    end
    always @(posedge \clk ) begin
        s582_val_n2 <= s581_val_n2;
    end
    always @(posedge \clk ) begin
        s582_val_n3 <= s581_val_n3;
    end
    always @(posedge \clk ) begin
        s582_val_n4 <= s581_val_n4;
    end
    always @(posedge \clk ) begin
        s582_val_n5 <= s581_val_n5;
    end
    always @(posedge \clk ) begin
        \s583_val  <= \s582_val ;
    end
    always @(posedge \clk ) begin
        s583_val_n1 <= s582_val_n1;
    end
    always @(posedge \clk ) begin
        s583_val_n2 <= s582_val_n2;
    end
    always @(posedge \clk ) begin
        s583_val_n3 <= s582_val_n3;
    end
    always @(posedge \clk ) begin
        s583_val_n4 <= s582_val_n4;
    end
    always @(posedge \clk ) begin
        s583_val_n5 <= s582_val_n5;
    end
    always @(posedge \clk ) begin
        \s584_val  <= \s583_val ;
    end
    always @(posedge \clk ) begin
        s584_val_n1 <= s583_val_n1;
    end
    always @(posedge \clk ) begin
        s584_val_n2 <= s583_val_n2;
    end
    always @(posedge \clk ) begin
        s584_val_n3 <= s583_val_n3;
    end
    always @(posedge \clk ) begin
        s584_val_n4 <= s583_val_n4;
    end
    always @(posedge \clk ) begin
        s584_val_n5 <= s583_val_n5;
    end
    always @(posedge \clk ) begin
        \s585_val  <= \s584_val ;
    end
    always @(posedge \clk ) begin
        s585_val_n1 <= s584_val_n1;
    end
    always @(posedge \clk ) begin
        s585_val_n2 <= s584_val_n2;
    end
    always @(posedge \clk ) begin
        s585_val_n3 <= s584_val_n3;
    end
    always @(posedge \clk ) begin
        s585_val_n4 <= s584_val_n4;
    end
    always @(posedge \clk ) begin
        s585_val_n5 <= s584_val_n5;
    end
    always @(posedge \clk ) begin
        \s586_val  <= \s585_val ;
    end
    always @(posedge \clk ) begin
        s586_val_n1 <= s585_val_n1;
    end
    always @(posedge \clk ) begin
        s586_val_n2 <= s585_val_n2;
    end
    always @(posedge \clk ) begin
        s586_val_n3 <= s585_val_n3;
    end
    always @(posedge \clk ) begin
        s586_val_n4 <= s585_val_n4;
    end
    always @(posedge \clk ) begin
        s586_val_n5 <= s585_val_n5;
    end
    always @(posedge \clk ) begin
        \s587_val  <= \s586_val ;
    end
    always @(posedge \clk ) begin
        s587_val_n1 <= s586_val_n1;
    end
    always @(posedge \clk ) begin
        s587_val_n2 <= s586_val_n2;
    end
    always @(posedge \clk ) begin
        s587_val_n3 <= s586_val_n3;
    end
    always @(posedge \clk ) begin
        s587_val_n4 <= s586_val_n4;
    end
    always @(posedge \clk ) begin
        s587_val_n5 <= s586_val_n5;
    end
    always @(posedge \clk ) begin
        \s588_val  <= \s587_val ;
    end
    always @(posedge \clk ) begin
        s588_val_n1 <= s587_val_n1;
    end
    always @(posedge \clk ) begin
        s588_val_n2 <= s587_val_n2;
    end
    always @(posedge \clk ) begin
        s588_val_n3 <= s587_val_n3;
    end
    always @(posedge \clk ) begin
        s588_val_n4 <= s587_val_n4;
    end
    always @(posedge \clk ) begin
        s588_val_n5 <= s587_val_n5;
    end
    always @(posedge \clk ) begin
        \s589_val  <= \s588_val ;
    end
    always @(posedge \clk ) begin
        s589_val_n1 <= s588_val_n1;
    end
    always @(posedge \clk ) begin
        s589_val_n2 <= s588_val_n2;
    end
    always @(posedge \clk ) begin
        s589_val_n3 <= s588_val_n3;
    end
    always @(posedge \clk ) begin
        s589_val_n4 <= s588_val_n4;
    end
    always @(posedge \clk ) begin
        s589_val_n5 <= s588_val_n5;
    end
    always @(posedge \clk ) begin
        \s590_val  <= \s589_val ;
    end
    always @(posedge \clk ) begin
        s590_val_n1 <= s589_val_n1;
    end
    always @(posedge \clk ) begin
        s590_val_n2 <= s589_val_n2;
    end
    always @(posedge \clk ) begin
        s590_val_n3 <= s589_val_n3;
    end
    always @(posedge \clk ) begin
        s590_val_n4 <= s589_val_n4;
    end
    always @(posedge \clk ) begin
        s590_val_n5 <= s589_val_n5;
    end
    always @(posedge \clk ) begin
        \s591_val  <= \s590_val ;
    end
    always @(posedge \clk ) begin
        s591_val_n1 <= s590_val_n1;
    end
    always @(posedge \clk ) begin
        s591_val_n2 <= s590_val_n2;
    end
    always @(posedge \clk ) begin
        s591_val_n3 <= s590_val_n3;
    end
    always @(posedge \clk ) begin
        s591_val_n4 <= s590_val_n4;
    end
    always @(posedge \clk ) begin
        s591_val_n5 <= s590_val_n5;
    end
    always @(posedge \clk ) begin
        \s592_val  <= \s591_val ;
    end
    always @(posedge \clk ) begin
        s592_val_n1 <= s591_val_n1;
    end
    always @(posedge \clk ) begin
        s592_val_n2 <= s591_val_n2;
    end
    always @(posedge \clk ) begin
        s592_val_n3 <= s591_val_n3;
    end
    always @(posedge \clk ) begin
        s592_val_n4 <= s591_val_n4;
    end
    always @(posedge \clk ) begin
        s592_val_n5 <= s591_val_n5;
    end
    always @(posedge \clk ) begin
        \s593_val  <= \s592_val ;
    end
    always @(posedge \clk ) begin
        s593_val_n1 <= s592_val_n1;
    end
    always @(posedge \clk ) begin
        s593_val_n2 <= s592_val_n2;
    end
    always @(posedge \clk ) begin
        s593_val_n3 <= s592_val_n3;
    end
    always @(posedge \clk ) begin
        s593_val_n4 <= s592_val_n4;
    end
    always @(posedge \clk ) begin
        s593_val_n5 <= s592_val_n5;
    end
    always @(posedge \clk ) begin
        \s594_val  <= \s593_val ;
    end
    always @(posedge \clk ) begin
        s594_val_n1 <= s593_val_n1;
    end
    always @(posedge \clk ) begin
        s594_val_n2 <= s593_val_n2;
    end
    always @(posedge \clk ) begin
        s594_val_n3 <= s593_val_n3;
    end
    always @(posedge \clk ) begin
        s594_val_n4 <= s593_val_n4;
    end
    always @(posedge \clk ) begin
        s594_val_n5 <= s593_val_n5;
    end
    always @(posedge \clk ) begin
        \s595_val  <= \s594_val ;
    end
    always @(posedge \clk ) begin
        s595_val_n1 <= s594_val_n1;
    end
    always @(posedge \clk ) begin
        s595_val_n2 <= s594_val_n2;
    end
    always @(posedge \clk ) begin
        s595_val_n3 <= s594_val_n3;
    end
    always @(posedge \clk ) begin
        s595_val_n4 <= s594_val_n4;
    end
    always @(posedge \clk ) begin
        s595_val_n5 <= s594_val_n5;
    end
    always @(posedge \clk ) begin
        \s596_val  <= \s595_val ;
    end
    always @(posedge \clk ) begin
        s596_val_n1 <= s595_val_n1;
    end
    always @(posedge \clk ) begin
        s596_val_n2 <= s595_val_n2;
    end
    always @(posedge \clk ) begin
        s596_val_n3 <= s595_val_n3;
    end
    always @(posedge \clk ) begin
        s596_val_n4 <= s595_val_n4;
    end
    always @(posedge \clk ) begin
        s596_val_n5 <= s595_val_n5;
    end
    always @(posedge \clk ) begin
        \s597_val  <= \s596_val ;
    end
    always @(posedge \clk ) begin
        s597_val_n1 <= s596_val_n1;
    end
    always @(posedge \clk ) begin
        s597_val_n2 <= s596_val_n2;
    end
    always @(posedge \clk ) begin
        s597_val_n3 <= s596_val_n3;
    end
    always @(posedge \clk ) begin
        s597_val_n4 <= s596_val_n4;
    end
    always @(posedge \clk ) begin
        s597_val_n5 <= s596_val_n5;
    end
    always @(posedge \clk ) begin
        \s598_val  <= \s597_val ;
    end
    always @(posedge \clk ) begin
        s598_val_n1 <= s597_val_n1;
    end
    always @(posedge \clk ) begin
        s598_val_n2 <= s597_val_n2;
    end
    always @(posedge \clk ) begin
        s598_val_n3 <= s597_val_n3;
    end
    always @(posedge \clk ) begin
        s598_val_n4 <= s597_val_n4;
    end
    always @(posedge \clk ) begin
        s598_val_n5 <= s597_val_n5;
    end
    always @(posedge \clk ) begin
        \s599_val  <= \s598_val ;
    end
    always @(posedge \clk ) begin
        s599_val_n1 <= s598_val_n1;
    end
    always @(posedge \clk ) begin
        s599_val_n2 <= s598_val_n2;
    end
    always @(posedge \clk ) begin
        s599_val_n3 <= s598_val_n3;
    end
    always @(posedge \clk ) begin
        s599_val_n4 <= s598_val_n4;
    end
    always @(posedge \clk ) begin
        s599_val_n5 <= s598_val_n5;
    end
    always @(posedge \clk ) begin
        \s600_val  <= \s599_val ;
    end
    always @(posedge \clk ) begin
        s600_val_n1 <= s599_val_n1;
    end
    always @(posedge \clk ) begin
        s600_val_n2 <= s599_val_n2;
    end
    always @(posedge \clk ) begin
        s600_val_n3 <= s599_val_n3;
    end
    always @(posedge \clk ) begin
        s600_val_n4 <= s599_val_n4;
    end
    always @(posedge \clk ) begin
        s600_val_n5 <= s599_val_n5;
    end
    always @(posedge \clk ) begin
        \s601_val  <= \s600_val ;
    end
    always @(posedge \clk ) begin
        s601_val_n1 <= s600_val_n1;
    end
    always @(posedge \clk ) begin
        s601_val_n2 <= s600_val_n2;
    end
    always @(posedge \clk ) begin
        s601_val_n3 <= s600_val_n3;
    end
    always @(posedge \clk ) begin
        s601_val_n4 <= s600_val_n4;
    end
    always @(posedge \clk ) begin
        s601_val_n5 <= s600_val_n5;
    end
    always @(posedge \clk ) begin
        s601_val_n6 <= val_n6;
    end
    always @(posedge \clk ) begin
        \s602_val  <= \s601_val ;
    end
    always @(posedge \clk ) begin
        s602_val_n1 <= s601_val_n1;
    end
    always @(posedge \clk ) begin
        s602_val_n2 <= s601_val_n2;
    end
    always @(posedge \clk ) begin
        s602_val_n3 <= s601_val_n3;
    end
    always @(posedge \clk ) begin
        s602_val_n4 <= s601_val_n4;
    end
    always @(posedge \clk ) begin
        s602_val_n5 <= s601_val_n5;
    end
    always @(posedge \clk ) begin
        s602_val_n6 <= s601_val_n6;
    end
    always @(posedge \clk ) begin
        \s603_val  <= \s602_val ;
    end
    always @(posedge \clk ) begin
        s603_val_n1 <= s602_val_n1;
    end
    always @(posedge \clk ) begin
        s603_val_n2 <= s602_val_n2;
    end
    always @(posedge \clk ) begin
        s603_val_n3 <= s602_val_n3;
    end
    always @(posedge \clk ) begin
        s603_val_n4 <= s602_val_n4;
    end
    always @(posedge \clk ) begin
        s603_val_n5 <= s602_val_n5;
    end
    always @(posedge \clk ) begin
        s603_val_n6 <= s602_val_n6;
    end
    always @(posedge \clk ) begin
        \s604_val  <= \s603_val ;
    end
    always @(posedge \clk ) begin
        s604_val_n1 <= s603_val_n1;
    end
    always @(posedge \clk ) begin
        s604_val_n2 <= s603_val_n2;
    end
    always @(posedge \clk ) begin
        s604_val_n3 <= s603_val_n3;
    end
    always @(posedge \clk ) begin
        s604_val_n4 <= s603_val_n4;
    end
    always @(posedge \clk ) begin
        s604_val_n5 <= s603_val_n5;
    end
    always @(posedge \clk ) begin
        s604_val_n6 <= s603_val_n6;
    end
    always @(posedge \clk ) begin
        \s605_val  <= \s604_val ;
    end
    always @(posedge \clk ) begin
        s605_val_n1 <= s604_val_n1;
    end
    always @(posedge \clk ) begin
        s605_val_n2 <= s604_val_n2;
    end
    always @(posedge \clk ) begin
        s605_val_n3 <= s604_val_n3;
    end
    always @(posedge \clk ) begin
        s605_val_n4 <= s604_val_n4;
    end
    always @(posedge \clk ) begin
        s605_val_n5 <= s604_val_n5;
    end
    always @(posedge \clk ) begin
        s605_val_n6 <= s604_val_n6;
    end
    always @(posedge \clk ) begin
        \s606_val  <= \s605_val ;
    end
    always @(posedge \clk ) begin
        s606_val_n1 <= s605_val_n1;
    end
    always @(posedge \clk ) begin
        s606_val_n2 <= s605_val_n2;
    end
    always @(posedge \clk ) begin
        s606_val_n3 <= s605_val_n3;
    end
    always @(posedge \clk ) begin
        s606_val_n4 <= s605_val_n4;
    end
    always @(posedge \clk ) begin
        s606_val_n5 <= s605_val_n5;
    end
    always @(posedge \clk ) begin
        s606_val_n6 <= s605_val_n6;
    end
    always @(posedge \clk ) begin
        \s607_val  <= \s606_val ;
    end
    always @(posedge \clk ) begin
        s607_val_n1 <= s606_val_n1;
    end
    always @(posedge \clk ) begin
        s607_val_n2 <= s606_val_n2;
    end
    always @(posedge \clk ) begin
        s607_val_n3 <= s606_val_n3;
    end
    always @(posedge \clk ) begin
        s607_val_n4 <= s606_val_n4;
    end
    always @(posedge \clk ) begin
        s607_val_n5 <= s606_val_n5;
    end
    always @(posedge \clk ) begin
        s607_val_n6 <= s606_val_n6;
    end
    always @(posedge \clk ) begin
        \s608_val  <= \s607_val ;
    end
    always @(posedge \clk ) begin
        s608_val_n1 <= s607_val_n1;
    end
    always @(posedge \clk ) begin
        s608_val_n2 <= s607_val_n2;
    end
    always @(posedge \clk ) begin
        s608_val_n3 <= s607_val_n3;
    end
    always @(posedge \clk ) begin
        s608_val_n4 <= s607_val_n4;
    end
    always @(posedge \clk ) begin
        s608_val_n5 <= s607_val_n5;
    end
    always @(posedge \clk ) begin
        s608_val_n6 <= s607_val_n6;
    end
    always @(posedge \clk ) begin
        \s609_val  <= \s608_val ;
    end
    always @(posedge \clk ) begin
        s609_val_n1 <= s608_val_n1;
    end
    always @(posedge \clk ) begin
        s609_val_n2 <= s608_val_n2;
    end
    always @(posedge \clk ) begin
        s609_val_n3 <= s608_val_n3;
    end
    always @(posedge \clk ) begin
        s609_val_n4 <= s608_val_n4;
    end
    always @(posedge \clk ) begin
        s609_val_n5 <= s608_val_n5;
    end
    always @(posedge \clk ) begin
        s609_val_n6 <= s608_val_n6;
    end
    always @(posedge \clk ) begin
        \s610_val  <= \s609_val ;
    end
    always @(posedge \clk ) begin
        s610_val_n1 <= s609_val_n1;
    end
    always @(posedge \clk ) begin
        s610_val_n2 <= s609_val_n2;
    end
    always @(posedge \clk ) begin
        s610_val_n3 <= s609_val_n3;
    end
    always @(posedge \clk ) begin
        s610_val_n4 <= s609_val_n4;
    end
    always @(posedge \clk ) begin
        s610_val_n5 <= s609_val_n5;
    end
    always @(posedge \clk ) begin
        s610_val_n6 <= s609_val_n6;
    end
    always @(posedge \clk ) begin
        \s611_val  <= \s610_val ;
    end
    always @(posedge \clk ) begin
        s611_val_n1 <= s610_val_n1;
    end
    always @(posedge \clk ) begin
        s611_val_n2 <= s610_val_n2;
    end
    always @(posedge \clk ) begin
        s611_val_n3 <= s610_val_n3;
    end
    always @(posedge \clk ) begin
        s611_val_n4 <= s610_val_n4;
    end
    always @(posedge \clk ) begin
        s611_val_n5 <= s610_val_n5;
    end
    always @(posedge \clk ) begin
        s611_val_n6 <= s610_val_n6;
    end
    always @(posedge \clk ) begin
        \s612_val  <= \s611_val ;
    end
    always @(posedge \clk ) begin
        s612_val_n1 <= s611_val_n1;
    end
    always @(posedge \clk ) begin
        s612_val_n2 <= s611_val_n2;
    end
    always @(posedge \clk ) begin
        s612_val_n3 <= s611_val_n3;
    end
    always @(posedge \clk ) begin
        s612_val_n4 <= s611_val_n4;
    end
    always @(posedge \clk ) begin
        s612_val_n5 <= s611_val_n5;
    end
    always @(posedge \clk ) begin
        s612_val_n6 <= s611_val_n6;
    end
    always @(posedge \clk ) begin
        \s613_val  <= \s612_val ;
    end
    always @(posedge \clk ) begin
        s613_val_n1 <= s612_val_n1;
    end
    always @(posedge \clk ) begin
        s613_val_n2 <= s612_val_n2;
    end
    always @(posedge \clk ) begin
        s613_val_n3 <= s612_val_n3;
    end
    always @(posedge \clk ) begin
        s613_val_n4 <= s612_val_n4;
    end
    always @(posedge \clk ) begin
        s613_val_n5 <= s612_val_n5;
    end
    always @(posedge \clk ) begin
        s613_val_n6 <= s612_val_n6;
    end
    always @(posedge \clk ) begin
        \s614_val  <= \s613_val ;
    end
    always @(posedge \clk ) begin
        s614_val_n1 <= s613_val_n1;
    end
    always @(posedge \clk ) begin
        s614_val_n2 <= s613_val_n2;
    end
    always @(posedge \clk ) begin
        s614_val_n3 <= s613_val_n3;
    end
    always @(posedge \clk ) begin
        s614_val_n4 <= s613_val_n4;
    end
    always @(posedge \clk ) begin
        s614_val_n5 <= s613_val_n5;
    end
    always @(posedge \clk ) begin
        s614_val_n6 <= s613_val_n6;
    end
    always @(posedge \clk ) begin
        \s615_val  <= \s614_val ;
    end
    always @(posedge \clk ) begin
        s615_val_n1 <= s614_val_n1;
    end
    always @(posedge \clk ) begin
        s615_val_n2 <= s614_val_n2;
    end
    always @(posedge \clk ) begin
        s615_val_n3 <= s614_val_n3;
    end
    always @(posedge \clk ) begin
        s615_val_n4 <= s614_val_n4;
    end
    always @(posedge \clk ) begin
        s615_val_n5 <= s614_val_n5;
    end
    always @(posedge \clk ) begin
        s615_val_n6 <= s614_val_n6;
    end
    always @(posedge \clk ) begin
        \s616_val  <= \s615_val ;
    end
    always @(posedge \clk ) begin
        s616_val_n1 <= s615_val_n1;
    end
    always @(posedge \clk ) begin
        s616_val_n2 <= s615_val_n2;
    end
    always @(posedge \clk ) begin
        s616_val_n3 <= s615_val_n3;
    end
    always @(posedge \clk ) begin
        s616_val_n4 <= s615_val_n4;
    end
    always @(posedge \clk ) begin
        s616_val_n5 <= s615_val_n5;
    end
    always @(posedge \clk ) begin
        s616_val_n6 <= s615_val_n6;
    end
    always @(posedge \clk ) begin
        \s617_val  <= \s616_val ;
    end
    always @(posedge \clk ) begin
        s617_val_n1 <= s616_val_n1;
    end
    always @(posedge \clk ) begin
        s617_val_n2 <= s616_val_n2;
    end
    always @(posedge \clk ) begin
        s617_val_n3 <= s616_val_n3;
    end
    always @(posedge \clk ) begin
        s617_val_n4 <= s616_val_n4;
    end
    always @(posedge \clk ) begin
        s617_val_n5 <= s616_val_n5;
    end
    always @(posedge \clk ) begin
        s617_val_n6 <= s616_val_n6;
    end
    always @(posedge \clk ) begin
        \s618_val  <= \s617_val ;
    end
    always @(posedge \clk ) begin
        s618_val_n1 <= s617_val_n1;
    end
    always @(posedge \clk ) begin
        s618_val_n2 <= s617_val_n2;
    end
    always @(posedge \clk ) begin
        s618_val_n3 <= s617_val_n3;
    end
    always @(posedge \clk ) begin
        s618_val_n4 <= s617_val_n4;
    end
    always @(posedge \clk ) begin
        s618_val_n5 <= s617_val_n5;
    end
    always @(posedge \clk ) begin
        s618_val_n6 <= s617_val_n6;
    end
    always @(posedge \clk ) begin
        \s619_val  <= \s618_val ;
    end
    always @(posedge \clk ) begin
        s619_val_n1 <= s618_val_n1;
    end
    always @(posedge \clk ) begin
        s619_val_n2 <= s618_val_n2;
    end
    always @(posedge \clk ) begin
        s619_val_n3 <= s618_val_n3;
    end
    always @(posedge \clk ) begin
        s619_val_n4 <= s618_val_n4;
    end
    always @(posedge \clk ) begin
        s619_val_n5 <= s618_val_n5;
    end
    always @(posedge \clk ) begin
        s619_val_n6 <= s618_val_n6;
    end
    always @(posedge \clk ) begin
        \s620_val  <= \s619_val ;
    end
    always @(posedge \clk ) begin
        s620_val_n1 <= s619_val_n1;
    end
    always @(posedge \clk ) begin
        s620_val_n2 <= s619_val_n2;
    end
    always @(posedge \clk ) begin
        s620_val_n3 <= s619_val_n3;
    end
    always @(posedge \clk ) begin
        s620_val_n4 <= s619_val_n4;
    end
    always @(posedge \clk ) begin
        s620_val_n5 <= s619_val_n5;
    end
    always @(posedge \clk ) begin
        s620_val_n6 <= s619_val_n6;
    end
    always @(posedge \clk ) begin
        \s621_val  <= \s620_val ;
    end
    always @(posedge \clk ) begin
        s621_val_n1 <= s620_val_n1;
    end
    always @(posedge \clk ) begin
        s621_val_n2 <= s620_val_n2;
    end
    always @(posedge \clk ) begin
        s621_val_n3 <= s620_val_n3;
    end
    always @(posedge \clk ) begin
        s621_val_n4 <= s620_val_n4;
    end
    always @(posedge \clk ) begin
        s621_val_n5 <= s620_val_n5;
    end
    always @(posedge \clk ) begin
        s621_val_n6 <= s620_val_n6;
    end
    always @(posedge \clk ) begin
        \s622_val  <= \s621_val ;
    end
    always @(posedge \clk ) begin
        s622_val_n1 <= s621_val_n1;
    end
    always @(posedge \clk ) begin
        s622_val_n2 <= s621_val_n2;
    end
    always @(posedge \clk ) begin
        s622_val_n3 <= s621_val_n3;
    end
    always @(posedge \clk ) begin
        s622_val_n4 <= s621_val_n4;
    end
    always @(posedge \clk ) begin
        s622_val_n5 <= s621_val_n5;
    end
    always @(posedge \clk ) begin
        s622_val_n6 <= s621_val_n6;
    end
    always @(posedge \clk ) begin
        \s623_val  <= \s622_val ;
    end
    always @(posedge \clk ) begin
        s623_val_n1 <= s622_val_n1;
    end
    always @(posedge \clk ) begin
        s623_val_n2 <= s622_val_n2;
    end
    always @(posedge \clk ) begin
        s623_val_n3 <= s622_val_n3;
    end
    always @(posedge \clk ) begin
        s623_val_n4 <= s622_val_n4;
    end
    always @(posedge \clk ) begin
        s623_val_n5 <= s622_val_n5;
    end
    always @(posedge \clk ) begin
        s623_val_n6 <= s622_val_n6;
    end
    always @(posedge \clk ) begin
        \s624_val  <= \s623_val ;
    end
    always @(posedge \clk ) begin
        s624_val_n1 <= s623_val_n1;
    end
    always @(posedge \clk ) begin
        s624_val_n2 <= s623_val_n2;
    end
    always @(posedge \clk ) begin
        s624_val_n3 <= s623_val_n3;
    end
    always @(posedge \clk ) begin
        s624_val_n4 <= s623_val_n4;
    end
    always @(posedge \clk ) begin
        s624_val_n5 <= s623_val_n5;
    end
    always @(posedge \clk ) begin
        s624_val_n6 <= s623_val_n6;
    end
    always @(posedge \clk ) begin
        \s625_val  <= \s624_val ;
    end
    always @(posedge \clk ) begin
        s625_val_n1 <= s624_val_n1;
    end
    always @(posedge \clk ) begin
        s625_val_n2 <= s624_val_n2;
    end
    always @(posedge \clk ) begin
        s625_val_n3 <= s624_val_n3;
    end
    always @(posedge \clk ) begin
        s625_val_n4 <= s624_val_n4;
    end
    always @(posedge \clk ) begin
        s625_val_n5 <= s624_val_n5;
    end
    always @(posedge \clk ) begin
        s625_val_n6 <= s624_val_n6;
    end
    always @(posedge \clk ) begin
        \s626_val  <= \s625_val ;
    end
    always @(posedge \clk ) begin
        s626_val_n1 <= s625_val_n1;
    end
    always @(posedge \clk ) begin
        s626_val_n2 <= s625_val_n2;
    end
    always @(posedge \clk ) begin
        s626_val_n3 <= s625_val_n3;
    end
    always @(posedge \clk ) begin
        s626_val_n4 <= s625_val_n4;
    end
    always @(posedge \clk ) begin
        s626_val_n5 <= s625_val_n5;
    end
    always @(posedge \clk ) begin
        s626_val_n6 <= s625_val_n6;
    end
    always @(posedge \clk ) begin
        \s627_val  <= \s626_val ;
    end
    always @(posedge \clk ) begin
        s627_val_n1 <= s626_val_n1;
    end
    always @(posedge \clk ) begin
        s627_val_n2 <= s626_val_n2;
    end
    always @(posedge \clk ) begin
        s627_val_n3 <= s626_val_n3;
    end
    always @(posedge \clk ) begin
        s627_val_n4 <= s626_val_n4;
    end
    always @(posedge \clk ) begin
        s627_val_n5 <= s626_val_n5;
    end
    always @(posedge \clk ) begin
        s627_val_n6 <= s626_val_n6;
    end
    always @(posedge \clk ) begin
        \s628_val  <= \s627_val ;
    end
    always @(posedge \clk ) begin
        s628_val_n1 <= s627_val_n1;
    end
    always @(posedge \clk ) begin
        s628_val_n2 <= s627_val_n2;
    end
    always @(posedge \clk ) begin
        s628_val_n3 <= s627_val_n3;
    end
    always @(posedge \clk ) begin
        s628_val_n4 <= s627_val_n4;
    end
    always @(posedge \clk ) begin
        s628_val_n5 <= s627_val_n5;
    end
    always @(posedge \clk ) begin
        s628_val_n6 <= s627_val_n6;
    end
    always @(posedge \clk ) begin
        \s629_val  <= \s628_val ;
    end
    always @(posedge \clk ) begin
        s629_val_n1 <= s628_val_n1;
    end
    always @(posedge \clk ) begin
        s629_val_n2 <= s628_val_n2;
    end
    always @(posedge \clk ) begin
        s629_val_n3 <= s628_val_n3;
    end
    always @(posedge \clk ) begin
        s629_val_n4 <= s628_val_n4;
    end
    always @(posedge \clk ) begin
        s629_val_n5 <= s628_val_n5;
    end
    always @(posedge \clk ) begin
        s629_val_n6 <= s628_val_n6;
    end
    always @(posedge \clk ) begin
        \s630_val  <= \s629_val ;
    end
    always @(posedge \clk ) begin
        s630_val_n1 <= s629_val_n1;
    end
    always @(posedge \clk ) begin
        s630_val_n2 <= s629_val_n2;
    end
    always @(posedge \clk ) begin
        s630_val_n3 <= s629_val_n3;
    end
    always @(posedge \clk ) begin
        s630_val_n4 <= s629_val_n4;
    end
    always @(posedge \clk ) begin
        s630_val_n5 <= s629_val_n5;
    end
    always @(posedge \clk ) begin
        s630_val_n6 <= s629_val_n6;
    end
    always @(posedge \clk ) begin
        \s631_val  <= \s630_val ;
    end
    always @(posedge \clk ) begin
        s631_val_n1 <= s630_val_n1;
    end
    always @(posedge \clk ) begin
        s631_val_n2 <= s630_val_n2;
    end
    always @(posedge \clk ) begin
        s631_val_n3 <= s630_val_n3;
    end
    always @(posedge \clk ) begin
        s631_val_n4 <= s630_val_n4;
    end
    always @(posedge \clk ) begin
        s631_val_n5 <= s630_val_n5;
    end
    always @(posedge \clk ) begin
        s631_val_n6 <= s630_val_n6;
    end
    always @(posedge \clk ) begin
        \s632_val  <= \s631_val ;
    end
    always @(posedge \clk ) begin
        s632_val_n1 <= s631_val_n1;
    end
    always @(posedge \clk ) begin
        s632_val_n2 <= s631_val_n2;
    end
    always @(posedge \clk ) begin
        s632_val_n3 <= s631_val_n3;
    end
    always @(posedge \clk ) begin
        s632_val_n4 <= s631_val_n4;
    end
    always @(posedge \clk ) begin
        s632_val_n5 <= s631_val_n5;
    end
    always @(posedge \clk ) begin
        s632_val_n6 <= s631_val_n6;
    end
    always @(posedge \clk ) begin
        \s633_val  <= \s632_val ;
    end
    always @(posedge \clk ) begin
        s633_val_n1 <= s632_val_n1;
    end
    always @(posedge \clk ) begin
        s633_val_n2 <= s632_val_n2;
    end
    always @(posedge \clk ) begin
        s633_val_n3 <= s632_val_n3;
    end
    always @(posedge \clk ) begin
        s633_val_n4 <= s632_val_n4;
    end
    always @(posedge \clk ) begin
        s633_val_n5 <= s632_val_n5;
    end
    always @(posedge \clk ) begin
        s633_val_n6 <= s632_val_n6;
    end
    always @(posedge \clk ) begin
        \s634_val  <= \s633_val ;
    end
    always @(posedge \clk ) begin
        s634_val_n1 <= s633_val_n1;
    end
    always @(posedge \clk ) begin
        s634_val_n2 <= s633_val_n2;
    end
    always @(posedge \clk ) begin
        s634_val_n3 <= s633_val_n3;
    end
    always @(posedge \clk ) begin
        s634_val_n4 <= s633_val_n4;
    end
    always @(posedge \clk ) begin
        s634_val_n5 <= s633_val_n5;
    end
    always @(posedge \clk ) begin
        s634_val_n6 <= s633_val_n6;
    end
    always @(posedge \clk ) begin
        \s635_val  <= \s634_val ;
    end
    always @(posedge \clk ) begin
        s635_val_n1 <= s634_val_n1;
    end
    always @(posedge \clk ) begin
        s635_val_n2 <= s634_val_n2;
    end
    always @(posedge \clk ) begin
        s635_val_n3 <= s634_val_n3;
    end
    always @(posedge \clk ) begin
        s635_val_n4 <= s634_val_n4;
    end
    always @(posedge \clk ) begin
        s635_val_n5 <= s634_val_n5;
    end
    always @(posedge \clk ) begin
        s635_val_n6 <= s634_val_n6;
    end
    always @(posedge \clk ) begin
        \s636_val  <= \s635_val ;
    end
    always @(posedge \clk ) begin
        s636_val_n1 <= s635_val_n1;
    end
    always @(posedge \clk ) begin
        s636_val_n2 <= s635_val_n2;
    end
    always @(posedge \clk ) begin
        s636_val_n3 <= s635_val_n3;
    end
    always @(posedge \clk ) begin
        s636_val_n4 <= s635_val_n4;
    end
    always @(posedge \clk ) begin
        s636_val_n5 <= s635_val_n5;
    end
    always @(posedge \clk ) begin
        s636_val_n6 <= s635_val_n6;
    end
    always @(posedge \clk ) begin
        \s637_val  <= \s636_val ;
    end
    always @(posedge \clk ) begin
        s637_val_n1 <= s636_val_n1;
    end
    always @(posedge \clk ) begin
        s637_val_n2 <= s636_val_n2;
    end
    always @(posedge \clk ) begin
        s637_val_n3 <= s636_val_n3;
    end
    always @(posedge \clk ) begin
        s637_val_n4 <= s636_val_n4;
    end
    always @(posedge \clk ) begin
        s637_val_n5 <= s636_val_n5;
    end
    always @(posedge \clk ) begin
        s637_val_n6 <= s636_val_n6;
    end
    always @(posedge \clk ) begin
        \s638_val  <= \s637_val ;
    end
    always @(posedge \clk ) begin
        s638_val_n1 <= s637_val_n1;
    end
    always @(posedge \clk ) begin
        s638_val_n2 <= s637_val_n2;
    end
    always @(posedge \clk ) begin
        s638_val_n3 <= s637_val_n3;
    end
    always @(posedge \clk ) begin
        s638_val_n4 <= s637_val_n4;
    end
    always @(posedge \clk ) begin
        s638_val_n5 <= s637_val_n5;
    end
    always @(posedge \clk ) begin
        s638_val_n6 <= s637_val_n6;
    end
    always @(posedge \clk ) begin
        \s639_val  <= \s638_val ;
    end
    always @(posedge \clk ) begin
        s639_val_n1 <= s638_val_n1;
    end
    always @(posedge \clk ) begin
        s639_val_n2 <= s638_val_n2;
    end
    always @(posedge \clk ) begin
        s639_val_n3 <= s638_val_n3;
    end
    always @(posedge \clk ) begin
        s639_val_n4 <= s638_val_n4;
    end
    always @(posedge \clk ) begin
        s639_val_n5 <= s638_val_n5;
    end
    always @(posedge \clk ) begin
        s639_val_n6 <= s638_val_n6;
    end
    always @(posedge \clk ) begin
        \s640_val  <= \s639_val ;
    end
    always @(posedge \clk ) begin
        s640_val_n1 <= s639_val_n1;
    end
    always @(posedge \clk ) begin
        s640_val_n2 <= s639_val_n2;
    end
    always @(posedge \clk ) begin
        s640_val_n3 <= s639_val_n3;
    end
    always @(posedge \clk ) begin
        s640_val_n4 <= s639_val_n4;
    end
    always @(posedge \clk ) begin
        s640_val_n5 <= s639_val_n5;
    end
    always @(posedge \clk ) begin
        s640_val_n6 <= s639_val_n6;
    end
    always @(posedge \clk ) begin
        \s641_val  <= \s640_val ;
    end
    always @(posedge \clk ) begin
        s641_val_n1 <= s640_val_n1;
    end
    always @(posedge \clk ) begin
        s641_val_n2 <= s640_val_n2;
    end
    always @(posedge \clk ) begin
        s641_val_n3 <= s640_val_n3;
    end
    always @(posedge \clk ) begin
        s641_val_n4 <= s640_val_n4;
    end
    always @(posedge \clk ) begin
        s641_val_n5 <= s640_val_n5;
    end
    always @(posedge \clk ) begin
        s641_val_n6 <= s640_val_n6;
    end
    always @(posedge \clk ) begin
        \s642_val  <= \s641_val ;
    end
    always @(posedge \clk ) begin
        s642_val_n1 <= s641_val_n1;
    end
    always @(posedge \clk ) begin
        s642_val_n2 <= s641_val_n2;
    end
    always @(posedge \clk ) begin
        s642_val_n3 <= s641_val_n3;
    end
    always @(posedge \clk ) begin
        s642_val_n4 <= s641_val_n4;
    end
    always @(posedge \clk ) begin
        s642_val_n5 <= s641_val_n5;
    end
    always @(posedge \clk ) begin
        s642_val_n6 <= s641_val_n6;
    end
    always @(posedge \clk ) begin
        \s643_val  <= \s642_val ;
    end
    always @(posedge \clk ) begin
        s643_val_n1 <= s642_val_n1;
    end
    always @(posedge \clk ) begin
        s643_val_n2 <= s642_val_n2;
    end
    always @(posedge \clk ) begin
        s643_val_n3 <= s642_val_n3;
    end
    always @(posedge \clk ) begin
        s643_val_n4 <= s642_val_n4;
    end
    always @(posedge \clk ) begin
        s643_val_n5 <= s642_val_n5;
    end
    always @(posedge \clk ) begin
        s643_val_n6 <= s642_val_n6;
    end
    always @(posedge \clk ) begin
        \s644_val  <= \s643_val ;
    end
    always @(posedge \clk ) begin
        s644_val_n1 <= s643_val_n1;
    end
    always @(posedge \clk ) begin
        s644_val_n2 <= s643_val_n2;
    end
    always @(posedge \clk ) begin
        s644_val_n3 <= s643_val_n3;
    end
    always @(posedge \clk ) begin
        s644_val_n4 <= s643_val_n4;
    end
    always @(posedge \clk ) begin
        s644_val_n5 <= s643_val_n5;
    end
    always @(posedge \clk ) begin
        s644_val_n6 <= s643_val_n6;
    end
    always @(posedge \clk ) begin
        \s645_val  <= \s644_val ;
    end
    always @(posedge \clk ) begin
        s645_val_n1 <= s644_val_n1;
    end
    always @(posedge \clk ) begin
        s645_val_n2 <= s644_val_n2;
    end
    always @(posedge \clk ) begin
        s645_val_n3 <= s644_val_n3;
    end
    always @(posedge \clk ) begin
        s645_val_n4 <= s644_val_n4;
    end
    always @(posedge \clk ) begin
        s645_val_n5 <= s644_val_n5;
    end
    always @(posedge \clk ) begin
        s645_val_n6 <= s644_val_n6;
    end
    always @(posedge \clk ) begin
        \s646_val  <= \s645_val ;
    end
    always @(posedge \clk ) begin
        s646_val_n1 <= s645_val_n1;
    end
    always @(posedge \clk ) begin
        s646_val_n2 <= s645_val_n2;
    end
    always @(posedge \clk ) begin
        s646_val_n3 <= s645_val_n3;
    end
    always @(posedge \clk ) begin
        s646_val_n4 <= s645_val_n4;
    end
    always @(posedge \clk ) begin
        s646_val_n5 <= s645_val_n5;
    end
    always @(posedge \clk ) begin
        s646_val_n6 <= s645_val_n6;
    end
    always @(posedge \clk ) begin
        \s647_val  <= \s646_val ;
    end
    always @(posedge \clk ) begin
        s647_val_n1 <= s646_val_n1;
    end
    always @(posedge \clk ) begin
        s647_val_n2 <= s646_val_n2;
    end
    always @(posedge \clk ) begin
        s647_val_n3 <= s646_val_n3;
    end
    always @(posedge \clk ) begin
        s647_val_n4 <= s646_val_n4;
    end
    always @(posedge \clk ) begin
        s647_val_n5 <= s646_val_n5;
    end
    always @(posedge \clk ) begin
        s647_val_n6 <= s646_val_n6;
    end
    always @(posedge \clk ) begin
        \s648_val  <= \s647_val ;
    end
    always @(posedge \clk ) begin
        s648_val_n1 <= s647_val_n1;
    end
    always @(posedge \clk ) begin
        s648_val_n2 <= s647_val_n2;
    end
    always @(posedge \clk ) begin
        s648_val_n3 <= s647_val_n3;
    end
    always @(posedge \clk ) begin
        s648_val_n4 <= s647_val_n4;
    end
    always @(posedge \clk ) begin
        s648_val_n5 <= s647_val_n5;
    end
    always @(posedge \clk ) begin
        s648_val_n6 <= s647_val_n6;
    end
    always @(posedge \clk ) begin
        \s649_val  <= \s648_val ;
    end
    always @(posedge \clk ) begin
        s649_val_n1 <= s648_val_n1;
    end
    always @(posedge \clk ) begin
        s649_val_n2 <= s648_val_n2;
    end
    always @(posedge \clk ) begin
        s649_val_n3 <= s648_val_n3;
    end
    always @(posedge \clk ) begin
        s649_val_n4 <= s648_val_n4;
    end
    always @(posedge \clk ) begin
        s649_val_n5 <= s648_val_n5;
    end
    always @(posedge \clk ) begin
        s649_val_n6 <= s648_val_n6;
    end
    always @(posedge \clk ) begin
        \s650_val  <= \s649_val ;
    end
    always @(posedge \clk ) begin
        s650_val_n1 <= s649_val_n1;
    end
    always @(posedge \clk ) begin
        s650_val_n2 <= s649_val_n2;
    end
    always @(posedge \clk ) begin
        s650_val_n3 <= s649_val_n3;
    end
    always @(posedge \clk ) begin
        s650_val_n4 <= s649_val_n4;
    end
    always @(posedge \clk ) begin
        s650_val_n5 <= s649_val_n5;
    end
    always @(posedge \clk ) begin
        s650_val_n6 <= s649_val_n6;
    end
    always @(posedge \clk ) begin
        \s651_val  <= \s650_val ;
    end
    always @(posedge \clk ) begin
        s651_val_n1 <= s650_val_n1;
    end
    always @(posedge \clk ) begin
        s651_val_n2 <= s650_val_n2;
    end
    always @(posedge \clk ) begin
        s651_val_n3 <= s650_val_n3;
    end
    always @(posedge \clk ) begin
        s651_val_n4 <= s650_val_n4;
    end
    always @(posedge \clk ) begin
        s651_val_n5 <= s650_val_n5;
    end
    always @(posedge \clk ) begin
        s651_val_n6 <= s650_val_n6;
    end
    always @(posedge \clk ) begin
        \s652_val  <= \s651_val ;
    end
    always @(posedge \clk ) begin
        s652_val_n1 <= s651_val_n1;
    end
    always @(posedge \clk ) begin
        s652_val_n2 <= s651_val_n2;
    end
    always @(posedge \clk ) begin
        s652_val_n3 <= s651_val_n3;
    end
    always @(posedge \clk ) begin
        s652_val_n4 <= s651_val_n4;
    end
    always @(posedge \clk ) begin
        s652_val_n5 <= s651_val_n5;
    end
    always @(posedge \clk ) begin
        s652_val_n6 <= s651_val_n6;
    end
    always @(posedge \clk ) begin
        \s653_val  <= \s652_val ;
    end
    always @(posedge \clk ) begin
        s653_val_n1 <= s652_val_n1;
    end
    always @(posedge \clk ) begin
        s653_val_n2 <= s652_val_n2;
    end
    always @(posedge \clk ) begin
        s653_val_n3 <= s652_val_n3;
    end
    always @(posedge \clk ) begin
        s653_val_n4 <= s652_val_n4;
    end
    always @(posedge \clk ) begin
        s653_val_n5 <= s652_val_n5;
    end
    always @(posedge \clk ) begin
        s653_val_n6 <= s652_val_n6;
    end
    always @(posedge \clk ) begin
        \s654_val  <= \s653_val ;
    end
    always @(posedge \clk ) begin
        s654_val_n1 <= s653_val_n1;
    end
    always @(posedge \clk ) begin
        s654_val_n2 <= s653_val_n2;
    end
    always @(posedge \clk ) begin
        s654_val_n3 <= s653_val_n3;
    end
    always @(posedge \clk ) begin
        s654_val_n4 <= s653_val_n4;
    end
    always @(posedge \clk ) begin
        s654_val_n5 <= s653_val_n5;
    end
    always @(posedge \clk ) begin
        s654_val_n6 <= s653_val_n6;
    end
    always @(posedge \clk ) begin
        \s655_val  <= \s654_val ;
    end
    always @(posedge \clk ) begin
        s655_val_n1 <= s654_val_n1;
    end
    always @(posedge \clk ) begin
        s655_val_n2 <= s654_val_n2;
    end
    always @(posedge \clk ) begin
        s655_val_n3 <= s654_val_n3;
    end
    always @(posedge \clk ) begin
        s655_val_n4 <= s654_val_n4;
    end
    always @(posedge \clk ) begin
        s655_val_n5 <= s654_val_n5;
    end
    always @(posedge \clk ) begin
        s655_val_n6 <= s654_val_n6;
    end
    always @(posedge \clk ) begin
        \s656_val  <= \s655_val ;
    end
    always @(posedge \clk ) begin
        s656_val_n1 <= s655_val_n1;
    end
    always @(posedge \clk ) begin
        s656_val_n2 <= s655_val_n2;
    end
    always @(posedge \clk ) begin
        s656_val_n3 <= s655_val_n3;
    end
    always @(posedge \clk ) begin
        s656_val_n4 <= s655_val_n4;
    end
    always @(posedge \clk ) begin
        s656_val_n5 <= s655_val_n5;
    end
    always @(posedge \clk ) begin
        s656_val_n6 <= s655_val_n6;
    end
    always @(posedge \clk ) begin
        \s657_val  <= \s656_val ;
    end
    always @(posedge \clk ) begin
        s657_val_n1 <= s656_val_n1;
    end
    always @(posedge \clk ) begin
        s657_val_n2 <= s656_val_n2;
    end
    always @(posedge \clk ) begin
        s657_val_n3 <= s656_val_n3;
    end
    always @(posedge \clk ) begin
        s657_val_n4 <= s656_val_n4;
    end
    always @(posedge \clk ) begin
        s657_val_n5 <= s656_val_n5;
    end
    always @(posedge \clk ) begin
        s657_val_n6 <= s656_val_n6;
    end
    always @(posedge \clk ) begin
        \s658_val  <= \s657_val ;
    end
    always @(posedge \clk ) begin
        s658_val_n1 <= s657_val_n1;
    end
    always @(posedge \clk ) begin
        s658_val_n2 <= s657_val_n2;
    end
    always @(posedge \clk ) begin
        s658_val_n3 <= s657_val_n3;
    end
    always @(posedge \clk ) begin
        s658_val_n4 <= s657_val_n4;
    end
    always @(posedge \clk ) begin
        s658_val_n5 <= s657_val_n5;
    end
    always @(posedge \clk ) begin
        s658_val_n6 <= s657_val_n6;
    end
    always @(posedge \clk ) begin
        \s659_val  <= \s658_val ;
    end
    always @(posedge \clk ) begin
        s659_val_n1 <= s658_val_n1;
    end
    always @(posedge \clk ) begin
        s659_val_n2 <= s658_val_n2;
    end
    always @(posedge \clk ) begin
        s659_val_n3 <= s658_val_n3;
    end
    always @(posedge \clk ) begin
        s659_val_n4 <= s658_val_n4;
    end
    always @(posedge \clk ) begin
        s659_val_n5 <= s658_val_n5;
    end
    always @(posedge \clk ) begin
        s659_val_n6 <= s658_val_n6;
    end
    always @(posedge \clk ) begin
        \s660_val  <= \s659_val ;
    end
    always @(posedge \clk ) begin
        s660_val_n1 <= s659_val_n1;
    end
    always @(posedge \clk ) begin
        s660_val_n2 <= s659_val_n2;
    end
    always @(posedge \clk ) begin
        s660_val_n3 <= s659_val_n3;
    end
    always @(posedge \clk ) begin
        s660_val_n4 <= s659_val_n4;
    end
    always @(posedge \clk ) begin
        s660_val_n5 <= s659_val_n5;
    end
    always @(posedge \clk ) begin
        s660_val_n6 <= s659_val_n6;
    end
    always @(posedge \clk ) begin
        \s661_val  <= \s660_val ;
    end
    always @(posedge \clk ) begin
        s661_val_n1 <= s660_val_n1;
    end
    always @(posedge \clk ) begin
        s661_val_n2 <= s660_val_n2;
    end
    always @(posedge \clk ) begin
        s661_val_n3 <= s660_val_n3;
    end
    always @(posedge \clk ) begin
        s661_val_n4 <= s660_val_n4;
    end
    always @(posedge \clk ) begin
        s661_val_n5 <= s660_val_n5;
    end
    always @(posedge \clk ) begin
        s661_val_n6 <= s660_val_n6;
    end
    always @(posedge \clk ) begin
        \s662_val  <= \s661_val ;
    end
    always @(posedge \clk ) begin
        s662_val_n1 <= s661_val_n1;
    end
    always @(posedge \clk ) begin
        s662_val_n2 <= s661_val_n2;
    end
    always @(posedge \clk ) begin
        s662_val_n3 <= s661_val_n3;
    end
    always @(posedge \clk ) begin
        s662_val_n4 <= s661_val_n4;
    end
    always @(posedge \clk ) begin
        s662_val_n5 <= s661_val_n5;
    end
    always @(posedge \clk ) begin
        s662_val_n6 <= s661_val_n6;
    end
    always @(posedge \clk ) begin
        \s663_val  <= \s662_val ;
    end
    always @(posedge \clk ) begin
        s663_val_n1 <= s662_val_n1;
    end
    always @(posedge \clk ) begin
        s663_val_n2 <= s662_val_n2;
    end
    always @(posedge \clk ) begin
        s663_val_n3 <= s662_val_n3;
    end
    always @(posedge \clk ) begin
        s663_val_n4 <= s662_val_n4;
    end
    always @(posedge \clk ) begin
        s663_val_n5 <= s662_val_n5;
    end
    always @(posedge \clk ) begin
        s663_val_n6 <= s662_val_n6;
    end
    always @(posedge \clk ) begin
        \s664_val  <= \s663_val ;
    end
    always @(posedge \clk ) begin
        s664_val_n1 <= s663_val_n1;
    end
    always @(posedge \clk ) begin
        s664_val_n2 <= s663_val_n2;
    end
    always @(posedge \clk ) begin
        s664_val_n3 <= s663_val_n3;
    end
    always @(posedge \clk ) begin
        s664_val_n4 <= s663_val_n4;
    end
    always @(posedge \clk ) begin
        s664_val_n5 <= s663_val_n5;
    end
    always @(posedge \clk ) begin
        s664_val_n6 <= s663_val_n6;
    end
    always @(posedge \clk ) begin
        \s665_val  <= \s664_val ;
    end
    always @(posedge \clk ) begin
        s665_val_n1 <= s664_val_n1;
    end
    always @(posedge \clk ) begin
        s665_val_n2 <= s664_val_n2;
    end
    always @(posedge \clk ) begin
        s665_val_n3 <= s664_val_n3;
    end
    always @(posedge \clk ) begin
        s665_val_n4 <= s664_val_n4;
    end
    always @(posedge \clk ) begin
        s665_val_n5 <= s664_val_n5;
    end
    always @(posedge \clk ) begin
        s665_val_n6 <= s664_val_n6;
    end
    always @(posedge \clk ) begin
        \s666_val  <= \s665_val ;
    end
    always @(posedge \clk ) begin
        s666_val_n1 <= s665_val_n1;
    end
    always @(posedge \clk ) begin
        s666_val_n2 <= s665_val_n2;
    end
    always @(posedge \clk ) begin
        s666_val_n3 <= s665_val_n3;
    end
    always @(posedge \clk ) begin
        s666_val_n4 <= s665_val_n4;
    end
    always @(posedge \clk ) begin
        s666_val_n5 <= s665_val_n5;
    end
    always @(posedge \clk ) begin
        s666_val_n6 <= s665_val_n6;
    end
    always @(posedge \clk ) begin
        \s667_val  <= \s666_val ;
    end
    always @(posedge \clk ) begin
        s667_val_n1 <= s666_val_n1;
    end
    always @(posedge \clk ) begin
        s667_val_n2 <= s666_val_n2;
    end
    always @(posedge \clk ) begin
        s667_val_n3 <= s666_val_n3;
    end
    always @(posedge \clk ) begin
        s667_val_n4 <= s666_val_n4;
    end
    always @(posedge \clk ) begin
        s667_val_n5 <= s666_val_n5;
    end
    always @(posedge \clk ) begin
        s667_val_n6 <= s666_val_n6;
    end
    always @(posedge \clk ) begin
        \s668_val  <= \s667_val ;
    end
    always @(posedge \clk ) begin
        s668_val_n1 <= s667_val_n1;
    end
    always @(posedge \clk ) begin
        s668_val_n2 <= s667_val_n2;
    end
    always @(posedge \clk ) begin
        s668_val_n3 <= s667_val_n3;
    end
    always @(posedge \clk ) begin
        s668_val_n4 <= s667_val_n4;
    end
    always @(posedge \clk ) begin
        s668_val_n5 <= s667_val_n5;
    end
    always @(posedge \clk ) begin
        s668_val_n6 <= s667_val_n6;
    end
    always @(posedge \clk ) begin
        \s669_val  <= \s668_val ;
    end
    always @(posedge \clk ) begin
        s669_val_n1 <= s668_val_n1;
    end
    always @(posedge \clk ) begin
        s669_val_n2 <= s668_val_n2;
    end
    always @(posedge \clk ) begin
        s669_val_n3 <= s668_val_n3;
    end
    always @(posedge \clk ) begin
        s669_val_n4 <= s668_val_n4;
    end
    always @(posedge \clk ) begin
        s669_val_n5 <= s668_val_n5;
    end
    always @(posedge \clk ) begin
        s669_val_n6 <= s668_val_n6;
    end
    always @(posedge \clk ) begin
        \s670_val  <= \s669_val ;
    end
    always @(posedge \clk ) begin
        s670_val_n1 <= s669_val_n1;
    end
    always @(posedge \clk ) begin
        s670_val_n2 <= s669_val_n2;
    end
    always @(posedge \clk ) begin
        s670_val_n3 <= s669_val_n3;
    end
    always @(posedge \clk ) begin
        s670_val_n4 <= s669_val_n4;
    end
    always @(posedge \clk ) begin
        s670_val_n5 <= s669_val_n5;
    end
    always @(posedge \clk ) begin
        s670_val_n6 <= s669_val_n6;
    end
    always @(posedge \clk ) begin
        \s671_val  <= \s670_val ;
    end
    always @(posedge \clk ) begin
        s671_val_n1 <= s670_val_n1;
    end
    always @(posedge \clk ) begin
        s671_val_n2 <= s670_val_n2;
    end
    always @(posedge \clk ) begin
        s671_val_n3 <= s670_val_n3;
    end
    always @(posedge \clk ) begin
        s671_val_n4 <= s670_val_n4;
    end
    always @(posedge \clk ) begin
        s671_val_n5 <= s670_val_n5;
    end
    always @(posedge \clk ) begin
        s671_val_n6 <= s670_val_n6;
    end
    always @(posedge \clk ) begin
        \s672_val  <= \s671_val ;
    end
    always @(posedge \clk ) begin
        s672_val_n1 <= s671_val_n1;
    end
    always @(posedge \clk ) begin
        s672_val_n2 <= s671_val_n2;
    end
    always @(posedge \clk ) begin
        s672_val_n3 <= s671_val_n3;
    end
    always @(posedge \clk ) begin
        s672_val_n4 <= s671_val_n4;
    end
    always @(posedge \clk ) begin
        s672_val_n5 <= s671_val_n5;
    end
    always @(posedge \clk ) begin
        s672_val_n6 <= s671_val_n6;
    end
    always @(posedge \clk ) begin
        \s673_val  <= \s672_val ;
    end
    always @(posedge \clk ) begin
        s673_val_n1 <= s672_val_n1;
    end
    always @(posedge \clk ) begin
        s673_val_n2 <= s672_val_n2;
    end
    always @(posedge \clk ) begin
        s673_val_n3 <= s672_val_n3;
    end
    always @(posedge \clk ) begin
        s673_val_n4 <= s672_val_n4;
    end
    always @(posedge \clk ) begin
        s673_val_n5 <= s672_val_n5;
    end
    always @(posedge \clk ) begin
        s673_val_n6 <= s672_val_n6;
    end
    always @(posedge \clk ) begin
        \s674_val  <= \s673_val ;
    end
    always @(posedge \clk ) begin
        s674_val_n1 <= s673_val_n1;
    end
    always @(posedge \clk ) begin
        s674_val_n2 <= s673_val_n2;
    end
    always @(posedge \clk ) begin
        s674_val_n3 <= s673_val_n3;
    end
    always @(posedge \clk ) begin
        s674_val_n4 <= s673_val_n4;
    end
    always @(posedge \clk ) begin
        s674_val_n5 <= s673_val_n5;
    end
    always @(posedge \clk ) begin
        s674_val_n6 <= s673_val_n6;
    end
    always @(posedge \clk ) begin
        \s675_val  <= \s674_val ;
    end
    always @(posedge \clk ) begin
        s675_val_n1 <= s674_val_n1;
    end
    always @(posedge \clk ) begin
        s675_val_n2 <= s674_val_n2;
    end
    always @(posedge \clk ) begin
        s675_val_n3 <= s674_val_n3;
    end
    always @(posedge \clk ) begin
        s675_val_n4 <= s674_val_n4;
    end
    always @(posedge \clk ) begin
        s675_val_n5 <= s674_val_n5;
    end
    always @(posedge \clk ) begin
        s675_val_n6 <= s674_val_n6;
    end
    always @(posedge \clk ) begin
        \s676_val  <= \s675_val ;
    end
    always @(posedge \clk ) begin
        s676_val_n1 <= s675_val_n1;
    end
    always @(posedge \clk ) begin
        s676_val_n2 <= s675_val_n2;
    end
    always @(posedge \clk ) begin
        s676_val_n3 <= s675_val_n3;
    end
    always @(posedge \clk ) begin
        s676_val_n4 <= s675_val_n4;
    end
    always @(posedge \clk ) begin
        s676_val_n5 <= s675_val_n5;
    end
    always @(posedge \clk ) begin
        s676_val_n6 <= s675_val_n6;
    end
    always @(posedge \clk ) begin
        \s677_val  <= \s676_val ;
    end
    always @(posedge \clk ) begin
        s677_val_n1 <= s676_val_n1;
    end
    always @(posedge \clk ) begin
        s677_val_n2 <= s676_val_n2;
    end
    always @(posedge \clk ) begin
        s677_val_n3 <= s676_val_n3;
    end
    always @(posedge \clk ) begin
        s677_val_n4 <= s676_val_n4;
    end
    always @(posedge \clk ) begin
        s677_val_n5 <= s676_val_n5;
    end
    always @(posedge \clk ) begin
        s677_val_n6 <= s676_val_n6;
    end
    always @(posedge \clk ) begin
        \s678_val  <= \s677_val ;
    end
    always @(posedge \clk ) begin
        s678_val_n1 <= s677_val_n1;
    end
    always @(posedge \clk ) begin
        s678_val_n2 <= s677_val_n2;
    end
    always @(posedge \clk ) begin
        s678_val_n3 <= s677_val_n3;
    end
    always @(posedge \clk ) begin
        s678_val_n4 <= s677_val_n4;
    end
    always @(posedge \clk ) begin
        s678_val_n5 <= s677_val_n5;
    end
    always @(posedge \clk ) begin
        s678_val_n6 <= s677_val_n6;
    end
    always @(posedge \clk ) begin
        \s679_val  <= \s678_val ;
    end
    always @(posedge \clk ) begin
        s679_val_n1 <= s678_val_n1;
    end
    always @(posedge \clk ) begin
        s679_val_n2 <= s678_val_n2;
    end
    always @(posedge \clk ) begin
        s679_val_n3 <= s678_val_n3;
    end
    always @(posedge \clk ) begin
        s679_val_n4 <= s678_val_n4;
    end
    always @(posedge \clk ) begin
        s679_val_n5 <= s678_val_n5;
    end
    always @(posedge \clk ) begin
        s679_val_n6 <= s678_val_n6;
    end
    always @(posedge \clk ) begin
        \s680_val  <= \s679_val ;
    end
    always @(posedge \clk ) begin
        s680_val_n1 <= s679_val_n1;
    end
    always @(posedge \clk ) begin
        s680_val_n2 <= s679_val_n2;
    end
    always @(posedge \clk ) begin
        s680_val_n3 <= s679_val_n3;
    end
    always @(posedge \clk ) begin
        s680_val_n4 <= s679_val_n4;
    end
    always @(posedge \clk ) begin
        s680_val_n5 <= s679_val_n5;
    end
    always @(posedge \clk ) begin
        s680_val_n6 <= s679_val_n6;
    end
    always @(posedge \clk ) begin
        \s681_val  <= \s680_val ;
    end
    always @(posedge \clk ) begin
        s681_val_n1 <= s680_val_n1;
    end
    always @(posedge \clk ) begin
        s681_val_n2 <= s680_val_n2;
    end
    always @(posedge \clk ) begin
        s681_val_n3 <= s680_val_n3;
    end
    always @(posedge \clk ) begin
        s681_val_n4 <= s680_val_n4;
    end
    always @(posedge \clk ) begin
        s681_val_n5 <= s680_val_n5;
    end
    always @(posedge \clk ) begin
        s681_val_n6 <= s680_val_n6;
    end
    always @(posedge \clk ) begin
        \s682_val  <= \s681_val ;
    end
    always @(posedge \clk ) begin
        s682_val_n1 <= s681_val_n1;
    end
    always @(posedge \clk ) begin
        s682_val_n2 <= s681_val_n2;
    end
    always @(posedge \clk ) begin
        s682_val_n3 <= s681_val_n3;
    end
    always @(posedge \clk ) begin
        s682_val_n4 <= s681_val_n4;
    end
    always @(posedge \clk ) begin
        s682_val_n5 <= s681_val_n5;
    end
    always @(posedge \clk ) begin
        s682_val_n6 <= s681_val_n6;
    end
    always @(posedge \clk ) begin
        \s683_val  <= \s682_val ;
    end
    always @(posedge \clk ) begin
        s683_val_n1 <= s682_val_n1;
    end
    always @(posedge \clk ) begin
        s683_val_n2 <= s682_val_n2;
    end
    always @(posedge \clk ) begin
        s683_val_n3 <= s682_val_n3;
    end
    always @(posedge \clk ) begin
        s683_val_n4 <= s682_val_n4;
    end
    always @(posedge \clk ) begin
        s683_val_n5 <= s682_val_n5;
    end
    always @(posedge \clk ) begin
        s683_val_n6 <= s682_val_n6;
    end
    always @(posedge \clk ) begin
        \s684_val  <= \s683_val ;
    end
    always @(posedge \clk ) begin
        s684_val_n1 <= s683_val_n1;
    end
    always @(posedge \clk ) begin
        s684_val_n2 <= s683_val_n2;
    end
    always @(posedge \clk ) begin
        s684_val_n3 <= s683_val_n3;
    end
    always @(posedge \clk ) begin
        s684_val_n4 <= s683_val_n4;
    end
    always @(posedge \clk ) begin
        s684_val_n5 <= s683_val_n5;
    end
    always @(posedge \clk ) begin
        s684_val_n6 <= s683_val_n6;
    end
    always @(posedge \clk ) begin
        \s685_val  <= \s684_val ;
    end
    always @(posedge \clk ) begin
        s685_val_n1 <= s684_val_n1;
    end
    always @(posedge \clk ) begin
        s685_val_n2 <= s684_val_n2;
    end
    always @(posedge \clk ) begin
        s685_val_n3 <= s684_val_n3;
    end
    always @(posedge \clk ) begin
        s685_val_n4 <= s684_val_n4;
    end
    always @(posedge \clk ) begin
        s685_val_n5 <= s684_val_n5;
    end
    always @(posedge \clk ) begin
        s685_val_n6 <= s684_val_n6;
    end
    always @(posedge \clk ) begin
        \s686_val  <= \s685_val ;
    end
    always @(posedge \clk ) begin
        s686_val_n1 <= s685_val_n1;
    end
    always @(posedge \clk ) begin
        s686_val_n2 <= s685_val_n2;
    end
    always @(posedge \clk ) begin
        s686_val_n3 <= s685_val_n3;
    end
    always @(posedge \clk ) begin
        s686_val_n4 <= s685_val_n4;
    end
    always @(posedge \clk ) begin
        s686_val_n5 <= s685_val_n5;
    end
    always @(posedge \clk ) begin
        s686_val_n6 <= s685_val_n6;
    end
    always @(posedge \clk ) begin
        \s687_val  <= \s686_val ;
    end
    always @(posedge \clk ) begin
        s687_val_n1 <= s686_val_n1;
    end
    always @(posedge \clk ) begin
        s687_val_n2 <= s686_val_n2;
    end
    always @(posedge \clk ) begin
        s687_val_n3 <= s686_val_n3;
    end
    always @(posedge \clk ) begin
        s687_val_n4 <= s686_val_n4;
    end
    always @(posedge \clk ) begin
        s687_val_n5 <= s686_val_n5;
    end
    always @(posedge \clk ) begin
        s687_val_n6 <= s686_val_n6;
    end
    always @(posedge \clk ) begin
        \s688_val  <= \s687_val ;
    end
    always @(posedge \clk ) begin
        s688_val_n1 <= s687_val_n1;
    end
    always @(posedge \clk ) begin
        s688_val_n2 <= s687_val_n2;
    end
    always @(posedge \clk ) begin
        s688_val_n3 <= s687_val_n3;
    end
    always @(posedge \clk ) begin
        s688_val_n4 <= s687_val_n4;
    end
    always @(posedge \clk ) begin
        s688_val_n5 <= s687_val_n5;
    end
    always @(posedge \clk ) begin
        s688_val_n6 <= s687_val_n6;
    end
    always @(posedge \clk ) begin
        \s689_val  <= \s688_val ;
    end
    always @(posedge \clk ) begin
        s689_val_n1 <= s688_val_n1;
    end
    always @(posedge \clk ) begin
        s689_val_n2 <= s688_val_n2;
    end
    always @(posedge \clk ) begin
        s689_val_n3 <= s688_val_n3;
    end
    always @(posedge \clk ) begin
        s689_val_n4 <= s688_val_n4;
    end
    always @(posedge \clk ) begin
        s689_val_n5 <= s688_val_n5;
    end
    always @(posedge \clk ) begin
        s689_val_n6 <= s688_val_n6;
    end
    always @(posedge \clk ) begin
        \s690_val  <= \s689_val ;
    end
    always @(posedge \clk ) begin
        s690_val_n1 <= s689_val_n1;
    end
    always @(posedge \clk ) begin
        s690_val_n2 <= s689_val_n2;
    end
    always @(posedge \clk ) begin
        s690_val_n3 <= s689_val_n3;
    end
    always @(posedge \clk ) begin
        s690_val_n4 <= s689_val_n4;
    end
    always @(posedge \clk ) begin
        s690_val_n5 <= s689_val_n5;
    end
    always @(posedge \clk ) begin
        s690_val_n6 <= s689_val_n6;
    end
    always @(posedge \clk ) begin
        \s691_val  <= \s690_val ;
    end
    always @(posedge \clk ) begin
        s691_val_n1 <= s690_val_n1;
    end
    always @(posedge \clk ) begin
        s691_val_n2 <= s690_val_n2;
    end
    always @(posedge \clk ) begin
        s691_val_n3 <= s690_val_n3;
    end
    always @(posedge \clk ) begin
        s691_val_n4 <= s690_val_n4;
    end
    always @(posedge \clk ) begin
        s691_val_n5 <= s690_val_n5;
    end
    always @(posedge \clk ) begin
        s691_val_n6 <= s690_val_n6;
    end
    always @(posedge \clk ) begin
        \s692_val  <= \s691_val ;
    end
    always @(posedge \clk ) begin
        s692_val_n1 <= s691_val_n1;
    end
    always @(posedge \clk ) begin
        s692_val_n2 <= s691_val_n2;
    end
    always @(posedge \clk ) begin
        s692_val_n3 <= s691_val_n3;
    end
    always @(posedge \clk ) begin
        s692_val_n4 <= s691_val_n4;
    end
    always @(posedge \clk ) begin
        s692_val_n5 <= s691_val_n5;
    end
    always @(posedge \clk ) begin
        s692_val_n6 <= s691_val_n6;
    end
    always @(posedge \clk ) begin
        \s693_val  <= \s692_val ;
    end
    always @(posedge \clk ) begin
        s693_val_n1 <= s692_val_n1;
    end
    always @(posedge \clk ) begin
        s693_val_n2 <= s692_val_n2;
    end
    always @(posedge \clk ) begin
        s693_val_n3 <= s692_val_n3;
    end
    always @(posedge \clk ) begin
        s693_val_n4 <= s692_val_n4;
    end
    always @(posedge \clk ) begin
        s693_val_n5 <= s692_val_n5;
    end
    always @(posedge \clk ) begin
        s693_val_n6 <= s692_val_n6;
    end
    always @(posedge \clk ) begin
        \s694_val  <= \s693_val ;
    end
    always @(posedge \clk ) begin
        s694_val_n1 <= s693_val_n1;
    end
    always @(posedge \clk ) begin
        s694_val_n2 <= s693_val_n2;
    end
    always @(posedge \clk ) begin
        s694_val_n3 <= s693_val_n3;
    end
    always @(posedge \clk ) begin
        s694_val_n4 <= s693_val_n4;
    end
    always @(posedge \clk ) begin
        s694_val_n5 <= s693_val_n5;
    end
    always @(posedge \clk ) begin
        s694_val_n6 <= s693_val_n6;
    end
    always @(posedge \clk ) begin
        \s695_val  <= \s694_val ;
    end
    always @(posedge \clk ) begin
        s695_val_n1 <= s694_val_n1;
    end
    always @(posedge \clk ) begin
        s695_val_n2 <= s694_val_n2;
    end
    always @(posedge \clk ) begin
        s695_val_n3 <= s694_val_n3;
    end
    always @(posedge \clk ) begin
        s695_val_n4 <= s694_val_n4;
    end
    always @(posedge \clk ) begin
        s695_val_n5 <= s694_val_n5;
    end
    always @(posedge \clk ) begin
        s695_val_n6 <= s694_val_n6;
    end
    always @(posedge \clk ) begin
        \s696_val  <= \s695_val ;
    end
    always @(posedge \clk ) begin
        s696_val_n1 <= s695_val_n1;
    end
    always @(posedge \clk ) begin
        s696_val_n2 <= s695_val_n2;
    end
    always @(posedge \clk ) begin
        s696_val_n3 <= s695_val_n3;
    end
    always @(posedge \clk ) begin
        s696_val_n4 <= s695_val_n4;
    end
    always @(posedge \clk ) begin
        s696_val_n5 <= s695_val_n5;
    end
    always @(posedge \clk ) begin
        s696_val_n6 <= s695_val_n6;
    end
    always @(posedge \clk ) begin
        \s697_val  <= \s696_val ;
    end
    always @(posedge \clk ) begin
        s697_val_n1 <= s696_val_n1;
    end
    always @(posedge \clk ) begin
        s697_val_n2 <= s696_val_n2;
    end
    always @(posedge \clk ) begin
        s697_val_n3 <= s696_val_n3;
    end
    always @(posedge \clk ) begin
        s697_val_n4 <= s696_val_n4;
    end
    always @(posedge \clk ) begin
        s697_val_n5 <= s696_val_n5;
    end
    always @(posedge \clk ) begin
        s697_val_n6 <= s696_val_n6;
    end
    always @(posedge \clk ) begin
        \s698_val  <= \s697_val ;
    end
    always @(posedge \clk ) begin
        s698_val_n1 <= s697_val_n1;
    end
    always @(posedge \clk ) begin
        s698_val_n2 <= s697_val_n2;
    end
    always @(posedge \clk ) begin
        s698_val_n3 <= s697_val_n3;
    end
    always @(posedge \clk ) begin
        s698_val_n4 <= s697_val_n4;
    end
    always @(posedge \clk ) begin
        s698_val_n5 <= s697_val_n5;
    end
    always @(posedge \clk ) begin
        s698_val_n6 <= s697_val_n6;
    end
    always @(posedge \clk ) begin
        \s699_val  <= \s698_val ;
    end
    always @(posedge \clk ) begin
        s699_val_n1 <= s698_val_n1;
    end
    always @(posedge \clk ) begin
        s699_val_n2 <= s698_val_n2;
    end
    always @(posedge \clk ) begin
        s699_val_n3 <= s698_val_n3;
    end
    always @(posedge \clk ) begin
        s699_val_n4 <= s698_val_n4;
    end
    always @(posedge \clk ) begin
        s699_val_n5 <= s698_val_n5;
    end
    always @(posedge \clk ) begin
        s699_val_n6 <= s698_val_n6;
    end
    always @(posedge \clk ) begin
        \s700_val  <= \s699_val ;
    end
    always @(posedge \clk ) begin
        s700_val_n1 <= s699_val_n1;
    end
    always @(posedge \clk ) begin
        s700_val_n2 <= s699_val_n2;
    end
    always @(posedge \clk ) begin
        s700_val_n3 <= s699_val_n3;
    end
    always @(posedge \clk ) begin
        s700_val_n4 <= s699_val_n4;
    end
    always @(posedge \clk ) begin
        s700_val_n5 <= s699_val_n5;
    end
    always @(posedge \clk ) begin
        s700_val_n6 <= s699_val_n6;
    end
    always @(posedge \clk ) begin
        \s701_val  <= \s700_val ;
    end
    always @(posedge \clk ) begin
        s701_val_n1 <= s700_val_n1;
    end
    always @(posedge \clk ) begin
        s701_val_n2 <= s700_val_n2;
    end
    always @(posedge \clk ) begin
        s701_val_n3 <= s700_val_n3;
    end
    always @(posedge \clk ) begin
        s701_val_n4 <= s700_val_n4;
    end
    always @(posedge \clk ) begin
        s701_val_n5 <= s700_val_n5;
    end
    always @(posedge \clk ) begin
        s701_val_n6 <= s700_val_n6;
    end
    always @(posedge \clk ) begin
        s701_val_n7 <= val_n7;
    end
    always @(posedge \clk ) begin
        \s702_val  <= \s701_val ;
    end
    always @(posedge \clk ) begin
        s702_val_n1 <= s701_val_n1;
    end
    always @(posedge \clk ) begin
        s702_val_n2 <= s701_val_n2;
    end
    always @(posedge \clk ) begin
        s702_val_n3 <= s701_val_n3;
    end
    always @(posedge \clk ) begin
        s702_val_n4 <= s701_val_n4;
    end
    always @(posedge \clk ) begin
        s702_val_n5 <= s701_val_n5;
    end
    always @(posedge \clk ) begin
        s702_val_n6 <= s701_val_n6;
    end
    always @(posedge \clk ) begin
        s702_val_n7 <= s701_val_n7;
    end
    always @(posedge \clk ) begin
        \s703_val  <= \s702_val ;
    end
    always @(posedge \clk ) begin
        s703_val_n1 <= s702_val_n1;
    end
    always @(posedge \clk ) begin
        s703_val_n2 <= s702_val_n2;
    end
    always @(posedge \clk ) begin
        s703_val_n3 <= s702_val_n3;
    end
    always @(posedge \clk ) begin
        s703_val_n4 <= s702_val_n4;
    end
    always @(posedge \clk ) begin
        s703_val_n5 <= s702_val_n5;
    end
    always @(posedge \clk ) begin
        s703_val_n6 <= s702_val_n6;
    end
    always @(posedge \clk ) begin
        s703_val_n7 <= s702_val_n7;
    end
    always @(posedge \clk ) begin
        \s704_val  <= \s703_val ;
    end
    always @(posedge \clk ) begin
        s704_val_n1 <= s703_val_n1;
    end
    always @(posedge \clk ) begin
        s704_val_n2 <= s703_val_n2;
    end
    always @(posedge \clk ) begin
        s704_val_n3 <= s703_val_n3;
    end
    always @(posedge \clk ) begin
        s704_val_n4 <= s703_val_n4;
    end
    always @(posedge \clk ) begin
        s704_val_n5 <= s703_val_n5;
    end
    always @(posedge \clk ) begin
        s704_val_n6 <= s703_val_n6;
    end
    always @(posedge \clk ) begin
        s704_val_n7 <= s703_val_n7;
    end
    always @(posedge \clk ) begin
        \s705_val  <= \s704_val ;
    end
    always @(posedge \clk ) begin
        s705_val_n1 <= s704_val_n1;
    end
    always @(posedge \clk ) begin
        s705_val_n2 <= s704_val_n2;
    end
    always @(posedge \clk ) begin
        s705_val_n3 <= s704_val_n3;
    end
    always @(posedge \clk ) begin
        s705_val_n4 <= s704_val_n4;
    end
    always @(posedge \clk ) begin
        s705_val_n5 <= s704_val_n5;
    end
    always @(posedge \clk ) begin
        s705_val_n6 <= s704_val_n6;
    end
    always @(posedge \clk ) begin
        s705_val_n7 <= s704_val_n7;
    end
    always @(posedge \clk ) begin
        \s706_val  <= \s705_val ;
    end
    always @(posedge \clk ) begin
        s706_val_n1 <= s705_val_n1;
    end
    always @(posedge \clk ) begin
        s706_val_n2 <= s705_val_n2;
    end
    always @(posedge \clk ) begin
        s706_val_n3 <= s705_val_n3;
    end
    always @(posedge \clk ) begin
        s706_val_n4 <= s705_val_n4;
    end
    always @(posedge \clk ) begin
        s706_val_n5 <= s705_val_n5;
    end
    always @(posedge \clk ) begin
        s706_val_n6 <= s705_val_n6;
    end
    always @(posedge \clk ) begin
        s706_val_n7 <= s705_val_n7;
    end
    always @(posedge \clk ) begin
        \s707_val  <= \s706_val ;
    end
    always @(posedge \clk ) begin
        s707_val_n1 <= s706_val_n1;
    end
    always @(posedge \clk ) begin
        s707_val_n2 <= s706_val_n2;
    end
    always @(posedge \clk ) begin
        s707_val_n3 <= s706_val_n3;
    end
    always @(posedge \clk ) begin
        s707_val_n4 <= s706_val_n4;
    end
    always @(posedge \clk ) begin
        s707_val_n5 <= s706_val_n5;
    end
    always @(posedge \clk ) begin
        s707_val_n6 <= s706_val_n6;
    end
    always @(posedge \clk ) begin
        s707_val_n7 <= s706_val_n7;
    end
    always @(posedge \clk ) begin
        \s708_val  <= \s707_val ;
    end
    always @(posedge \clk ) begin
        s708_val_n1 <= s707_val_n1;
    end
    always @(posedge \clk ) begin
        s708_val_n2 <= s707_val_n2;
    end
    always @(posedge \clk ) begin
        s708_val_n3 <= s707_val_n3;
    end
    always @(posedge \clk ) begin
        s708_val_n4 <= s707_val_n4;
    end
    always @(posedge \clk ) begin
        s708_val_n5 <= s707_val_n5;
    end
    always @(posedge \clk ) begin
        s708_val_n6 <= s707_val_n6;
    end
    always @(posedge \clk ) begin
        s708_val_n7 <= s707_val_n7;
    end
    always @(posedge \clk ) begin
        \s709_val  <= \s708_val ;
    end
    always @(posedge \clk ) begin
        s709_val_n1 <= s708_val_n1;
    end
    always @(posedge \clk ) begin
        s709_val_n2 <= s708_val_n2;
    end
    always @(posedge \clk ) begin
        s709_val_n3 <= s708_val_n3;
    end
    always @(posedge \clk ) begin
        s709_val_n4 <= s708_val_n4;
    end
    always @(posedge \clk ) begin
        s709_val_n5 <= s708_val_n5;
    end
    always @(posedge \clk ) begin
        s709_val_n6 <= s708_val_n6;
    end
    always @(posedge \clk ) begin
        s709_val_n7 <= s708_val_n7;
    end
    always @(posedge \clk ) begin
        \s710_val  <= \s709_val ;
    end
    always @(posedge \clk ) begin
        s710_val_n1 <= s709_val_n1;
    end
    always @(posedge \clk ) begin
        s710_val_n2 <= s709_val_n2;
    end
    always @(posedge \clk ) begin
        s710_val_n3 <= s709_val_n3;
    end
    always @(posedge \clk ) begin
        s710_val_n4 <= s709_val_n4;
    end
    always @(posedge \clk ) begin
        s710_val_n5 <= s709_val_n5;
    end
    always @(posedge \clk ) begin
        s710_val_n6 <= s709_val_n6;
    end
    always @(posedge \clk ) begin
        s710_val_n7 <= s709_val_n7;
    end
    always @(posedge \clk ) begin
        \s711_val  <= \s710_val ;
    end
    always @(posedge \clk ) begin
        s711_val_n1 <= s710_val_n1;
    end
    always @(posedge \clk ) begin
        s711_val_n2 <= s710_val_n2;
    end
    always @(posedge \clk ) begin
        s711_val_n3 <= s710_val_n3;
    end
    always @(posedge \clk ) begin
        s711_val_n4 <= s710_val_n4;
    end
    always @(posedge \clk ) begin
        s711_val_n5 <= s710_val_n5;
    end
    always @(posedge \clk ) begin
        s711_val_n6 <= s710_val_n6;
    end
    always @(posedge \clk ) begin
        s711_val_n7 <= s710_val_n7;
    end
    always @(posedge \clk ) begin
        \s712_val  <= \s711_val ;
    end
    always @(posedge \clk ) begin
        s712_val_n1 <= s711_val_n1;
    end
    always @(posedge \clk ) begin
        s712_val_n2 <= s711_val_n2;
    end
    always @(posedge \clk ) begin
        s712_val_n3 <= s711_val_n3;
    end
    always @(posedge \clk ) begin
        s712_val_n4 <= s711_val_n4;
    end
    always @(posedge \clk ) begin
        s712_val_n5 <= s711_val_n5;
    end
    always @(posedge \clk ) begin
        s712_val_n6 <= s711_val_n6;
    end
    always @(posedge \clk ) begin
        s712_val_n7 <= s711_val_n7;
    end
    always @(posedge \clk ) begin
        \s713_val  <= \s712_val ;
    end
    always @(posedge \clk ) begin
        s713_val_n1 <= s712_val_n1;
    end
    always @(posedge \clk ) begin
        s713_val_n2 <= s712_val_n2;
    end
    always @(posedge \clk ) begin
        s713_val_n3 <= s712_val_n3;
    end
    always @(posedge \clk ) begin
        s713_val_n4 <= s712_val_n4;
    end
    always @(posedge \clk ) begin
        s713_val_n5 <= s712_val_n5;
    end
    always @(posedge \clk ) begin
        s713_val_n6 <= s712_val_n6;
    end
    always @(posedge \clk ) begin
        s713_val_n7 <= s712_val_n7;
    end
    always @(posedge \clk ) begin
        \s714_val  <= \s713_val ;
    end
    always @(posedge \clk ) begin
        s714_val_n1 <= s713_val_n1;
    end
    always @(posedge \clk ) begin
        s714_val_n2 <= s713_val_n2;
    end
    always @(posedge \clk ) begin
        s714_val_n3 <= s713_val_n3;
    end
    always @(posedge \clk ) begin
        s714_val_n4 <= s713_val_n4;
    end
    always @(posedge \clk ) begin
        s714_val_n5 <= s713_val_n5;
    end
    always @(posedge \clk ) begin
        s714_val_n6 <= s713_val_n6;
    end
    always @(posedge \clk ) begin
        s714_val_n7 <= s713_val_n7;
    end
    always @(posedge \clk ) begin
        \s715_val  <= \s714_val ;
    end
    always @(posedge \clk ) begin
        s715_val_n1 <= s714_val_n1;
    end
    always @(posedge \clk ) begin
        s715_val_n2 <= s714_val_n2;
    end
    always @(posedge \clk ) begin
        s715_val_n3 <= s714_val_n3;
    end
    always @(posedge \clk ) begin
        s715_val_n4 <= s714_val_n4;
    end
    always @(posedge \clk ) begin
        s715_val_n5 <= s714_val_n5;
    end
    always @(posedge \clk ) begin
        s715_val_n6 <= s714_val_n6;
    end
    always @(posedge \clk ) begin
        s715_val_n7 <= s714_val_n7;
    end
    always @(posedge \clk ) begin
        \s716_val  <= \s715_val ;
    end
    always @(posedge \clk ) begin
        s716_val_n1 <= s715_val_n1;
    end
    always @(posedge \clk ) begin
        s716_val_n2 <= s715_val_n2;
    end
    always @(posedge \clk ) begin
        s716_val_n3 <= s715_val_n3;
    end
    always @(posedge \clk ) begin
        s716_val_n4 <= s715_val_n4;
    end
    always @(posedge \clk ) begin
        s716_val_n5 <= s715_val_n5;
    end
    always @(posedge \clk ) begin
        s716_val_n6 <= s715_val_n6;
    end
    always @(posedge \clk ) begin
        s716_val_n7 <= s715_val_n7;
    end
    always @(posedge \clk ) begin
        \s717_val  <= \s716_val ;
    end
    always @(posedge \clk ) begin
        s717_val_n1 <= s716_val_n1;
    end
    always @(posedge \clk ) begin
        s717_val_n2 <= s716_val_n2;
    end
    always @(posedge \clk ) begin
        s717_val_n3 <= s716_val_n3;
    end
    always @(posedge \clk ) begin
        s717_val_n4 <= s716_val_n4;
    end
    always @(posedge \clk ) begin
        s717_val_n5 <= s716_val_n5;
    end
    always @(posedge \clk ) begin
        s717_val_n6 <= s716_val_n6;
    end
    always @(posedge \clk ) begin
        s717_val_n7 <= s716_val_n7;
    end
    always @(posedge \clk ) begin
        \s718_val  <= \s717_val ;
    end
    always @(posedge \clk ) begin
        s718_val_n1 <= s717_val_n1;
    end
    always @(posedge \clk ) begin
        s718_val_n2 <= s717_val_n2;
    end
    always @(posedge \clk ) begin
        s718_val_n3 <= s717_val_n3;
    end
    always @(posedge \clk ) begin
        s718_val_n4 <= s717_val_n4;
    end
    always @(posedge \clk ) begin
        s718_val_n5 <= s717_val_n5;
    end
    always @(posedge \clk ) begin
        s718_val_n6 <= s717_val_n6;
    end
    always @(posedge \clk ) begin
        s718_val_n7 <= s717_val_n7;
    end
    always @(posedge \clk ) begin
        \s719_val  <= \s718_val ;
    end
    always @(posedge \clk ) begin
        s719_val_n1 <= s718_val_n1;
    end
    always @(posedge \clk ) begin
        s719_val_n2 <= s718_val_n2;
    end
    always @(posedge \clk ) begin
        s719_val_n3 <= s718_val_n3;
    end
    always @(posedge \clk ) begin
        s719_val_n4 <= s718_val_n4;
    end
    always @(posedge \clk ) begin
        s719_val_n5 <= s718_val_n5;
    end
    always @(posedge \clk ) begin
        s719_val_n6 <= s718_val_n6;
    end
    always @(posedge \clk ) begin
        s719_val_n7 <= s718_val_n7;
    end
    always @(posedge \clk ) begin
        \s720_val  <= \s719_val ;
    end
    always @(posedge \clk ) begin
        s720_val_n1 <= s719_val_n1;
    end
    always @(posedge \clk ) begin
        s720_val_n2 <= s719_val_n2;
    end
    always @(posedge \clk ) begin
        s720_val_n3 <= s719_val_n3;
    end
    always @(posedge \clk ) begin
        s720_val_n4 <= s719_val_n4;
    end
    always @(posedge \clk ) begin
        s720_val_n5 <= s719_val_n5;
    end
    always @(posedge \clk ) begin
        s720_val_n6 <= s719_val_n6;
    end
    always @(posedge \clk ) begin
        s720_val_n7 <= s719_val_n7;
    end
    always @(posedge \clk ) begin
        \s721_val  <= \s720_val ;
    end
    always @(posedge \clk ) begin
        s721_val_n1 <= s720_val_n1;
    end
    always @(posedge \clk ) begin
        s721_val_n2 <= s720_val_n2;
    end
    always @(posedge \clk ) begin
        s721_val_n3 <= s720_val_n3;
    end
    always @(posedge \clk ) begin
        s721_val_n4 <= s720_val_n4;
    end
    always @(posedge \clk ) begin
        s721_val_n5 <= s720_val_n5;
    end
    always @(posedge \clk ) begin
        s721_val_n6 <= s720_val_n6;
    end
    always @(posedge \clk ) begin
        s721_val_n7 <= s720_val_n7;
    end
    always @(posedge \clk ) begin
        \s722_val  <= \s721_val ;
    end
    always @(posedge \clk ) begin
        s722_val_n1 <= s721_val_n1;
    end
    always @(posedge \clk ) begin
        s722_val_n2 <= s721_val_n2;
    end
    always @(posedge \clk ) begin
        s722_val_n3 <= s721_val_n3;
    end
    always @(posedge \clk ) begin
        s722_val_n4 <= s721_val_n4;
    end
    always @(posedge \clk ) begin
        s722_val_n5 <= s721_val_n5;
    end
    always @(posedge \clk ) begin
        s722_val_n6 <= s721_val_n6;
    end
    always @(posedge \clk ) begin
        s722_val_n7 <= s721_val_n7;
    end
    always @(posedge \clk ) begin
        \s723_val  <= \s722_val ;
    end
    always @(posedge \clk ) begin
        s723_val_n1 <= s722_val_n1;
    end
    always @(posedge \clk ) begin
        s723_val_n2 <= s722_val_n2;
    end
    always @(posedge \clk ) begin
        s723_val_n3 <= s722_val_n3;
    end
    always @(posedge \clk ) begin
        s723_val_n4 <= s722_val_n4;
    end
    always @(posedge \clk ) begin
        s723_val_n5 <= s722_val_n5;
    end
    always @(posedge \clk ) begin
        s723_val_n6 <= s722_val_n6;
    end
    always @(posedge \clk ) begin
        s723_val_n7 <= s722_val_n7;
    end
    always @(posedge \clk ) begin
        \s724_val  <= \s723_val ;
    end
    always @(posedge \clk ) begin
        s724_val_n1 <= s723_val_n1;
    end
    always @(posedge \clk ) begin
        s724_val_n2 <= s723_val_n2;
    end
    always @(posedge \clk ) begin
        s724_val_n3 <= s723_val_n3;
    end
    always @(posedge \clk ) begin
        s724_val_n4 <= s723_val_n4;
    end
    always @(posedge \clk ) begin
        s724_val_n5 <= s723_val_n5;
    end
    always @(posedge \clk ) begin
        s724_val_n6 <= s723_val_n6;
    end
    always @(posedge \clk ) begin
        s724_val_n7 <= s723_val_n7;
    end
    always @(posedge \clk ) begin
        \s725_val  <= \s724_val ;
    end
    always @(posedge \clk ) begin
        s725_val_n1 <= s724_val_n1;
    end
    always @(posedge \clk ) begin
        s725_val_n2 <= s724_val_n2;
    end
    always @(posedge \clk ) begin
        s725_val_n3 <= s724_val_n3;
    end
    always @(posedge \clk ) begin
        s725_val_n4 <= s724_val_n4;
    end
    always @(posedge \clk ) begin
        s725_val_n5 <= s724_val_n5;
    end
    always @(posedge \clk ) begin
        s725_val_n6 <= s724_val_n6;
    end
    always @(posedge \clk ) begin
        s725_val_n7 <= s724_val_n7;
    end
    always @(posedge \clk ) begin
        \s726_val  <= \s725_val ;
    end
    always @(posedge \clk ) begin
        s726_val_n1 <= s725_val_n1;
    end
    always @(posedge \clk ) begin
        s726_val_n2 <= s725_val_n2;
    end
    always @(posedge \clk ) begin
        s726_val_n3 <= s725_val_n3;
    end
    always @(posedge \clk ) begin
        s726_val_n4 <= s725_val_n4;
    end
    always @(posedge \clk ) begin
        s726_val_n5 <= s725_val_n5;
    end
    always @(posedge \clk ) begin
        s726_val_n6 <= s725_val_n6;
    end
    always @(posedge \clk ) begin
        s726_val_n7 <= s725_val_n7;
    end
    always @(posedge \clk ) begin
        \s727_val  <= \s726_val ;
    end
    always @(posedge \clk ) begin
        s727_val_n1 <= s726_val_n1;
    end
    always @(posedge \clk ) begin
        s727_val_n2 <= s726_val_n2;
    end
    always @(posedge \clk ) begin
        s727_val_n3 <= s726_val_n3;
    end
    always @(posedge \clk ) begin
        s727_val_n4 <= s726_val_n4;
    end
    always @(posedge \clk ) begin
        s727_val_n5 <= s726_val_n5;
    end
    always @(posedge \clk ) begin
        s727_val_n6 <= s726_val_n6;
    end
    always @(posedge \clk ) begin
        s727_val_n7 <= s726_val_n7;
    end
    always @(posedge \clk ) begin
        \s728_val  <= \s727_val ;
    end
    always @(posedge \clk ) begin
        s728_val_n1 <= s727_val_n1;
    end
    always @(posedge \clk ) begin
        s728_val_n2 <= s727_val_n2;
    end
    always @(posedge \clk ) begin
        s728_val_n3 <= s727_val_n3;
    end
    always @(posedge \clk ) begin
        s728_val_n4 <= s727_val_n4;
    end
    always @(posedge \clk ) begin
        s728_val_n5 <= s727_val_n5;
    end
    always @(posedge \clk ) begin
        s728_val_n6 <= s727_val_n6;
    end
    always @(posedge \clk ) begin
        s728_val_n7 <= s727_val_n7;
    end
    always @(posedge \clk ) begin
        \s729_val  <= \s728_val ;
    end
    always @(posedge \clk ) begin
        s729_val_n1 <= s728_val_n1;
    end
    always @(posedge \clk ) begin
        s729_val_n2 <= s728_val_n2;
    end
    always @(posedge \clk ) begin
        s729_val_n3 <= s728_val_n3;
    end
    always @(posedge \clk ) begin
        s729_val_n4 <= s728_val_n4;
    end
    always @(posedge \clk ) begin
        s729_val_n5 <= s728_val_n5;
    end
    always @(posedge \clk ) begin
        s729_val_n6 <= s728_val_n6;
    end
    always @(posedge \clk ) begin
        s729_val_n7 <= s728_val_n7;
    end
    always @(posedge \clk ) begin
        \s730_val  <= \s729_val ;
    end
    always @(posedge \clk ) begin
        s730_val_n1 <= s729_val_n1;
    end
    always @(posedge \clk ) begin
        s730_val_n2 <= s729_val_n2;
    end
    always @(posedge \clk ) begin
        s730_val_n3 <= s729_val_n3;
    end
    always @(posedge \clk ) begin
        s730_val_n4 <= s729_val_n4;
    end
    always @(posedge \clk ) begin
        s730_val_n5 <= s729_val_n5;
    end
    always @(posedge \clk ) begin
        s730_val_n6 <= s729_val_n6;
    end
    always @(posedge \clk ) begin
        s730_val_n7 <= s729_val_n7;
    end
    always @(posedge \clk ) begin
        \s731_val  <= \s730_val ;
    end
    always @(posedge \clk ) begin
        s731_val_n1 <= s730_val_n1;
    end
    always @(posedge \clk ) begin
        s731_val_n2 <= s730_val_n2;
    end
    always @(posedge \clk ) begin
        s731_val_n3 <= s730_val_n3;
    end
    always @(posedge \clk ) begin
        s731_val_n4 <= s730_val_n4;
    end
    always @(posedge \clk ) begin
        s731_val_n5 <= s730_val_n5;
    end
    always @(posedge \clk ) begin
        s731_val_n6 <= s730_val_n6;
    end
    always @(posedge \clk ) begin
        s731_val_n7 <= s730_val_n7;
    end
    always @(posedge \clk ) begin
        \s732_val  <= \s731_val ;
    end
    always @(posedge \clk ) begin
        s732_val_n1 <= s731_val_n1;
    end
    always @(posedge \clk ) begin
        s732_val_n2 <= s731_val_n2;
    end
    always @(posedge \clk ) begin
        s732_val_n3 <= s731_val_n3;
    end
    always @(posedge \clk ) begin
        s732_val_n4 <= s731_val_n4;
    end
    always @(posedge \clk ) begin
        s732_val_n5 <= s731_val_n5;
    end
    always @(posedge \clk ) begin
        s732_val_n6 <= s731_val_n6;
    end
    always @(posedge \clk ) begin
        s732_val_n7 <= s731_val_n7;
    end
    always @(posedge \clk ) begin
        \s733_val  <= \s732_val ;
    end
    always @(posedge \clk ) begin
        s733_val_n1 <= s732_val_n1;
    end
    always @(posedge \clk ) begin
        s733_val_n2 <= s732_val_n2;
    end
    always @(posedge \clk ) begin
        s733_val_n3 <= s732_val_n3;
    end
    always @(posedge \clk ) begin
        s733_val_n4 <= s732_val_n4;
    end
    always @(posedge \clk ) begin
        s733_val_n5 <= s732_val_n5;
    end
    always @(posedge \clk ) begin
        s733_val_n6 <= s732_val_n6;
    end
    always @(posedge \clk ) begin
        s733_val_n7 <= s732_val_n7;
    end
    always @(posedge \clk ) begin
        \s734_val  <= \s733_val ;
    end
    always @(posedge \clk ) begin
        s734_val_n1 <= s733_val_n1;
    end
    always @(posedge \clk ) begin
        s734_val_n2 <= s733_val_n2;
    end
    always @(posedge \clk ) begin
        s734_val_n3 <= s733_val_n3;
    end
    always @(posedge \clk ) begin
        s734_val_n4 <= s733_val_n4;
    end
    always @(posedge \clk ) begin
        s734_val_n5 <= s733_val_n5;
    end
    always @(posedge \clk ) begin
        s734_val_n6 <= s733_val_n6;
    end
    always @(posedge \clk ) begin
        s734_val_n7 <= s733_val_n7;
    end
    always @(posedge \clk ) begin
        \s735_val  <= \s734_val ;
    end
    always @(posedge \clk ) begin
        s735_val_n1 <= s734_val_n1;
    end
    always @(posedge \clk ) begin
        s735_val_n2 <= s734_val_n2;
    end
    always @(posedge \clk ) begin
        s735_val_n3 <= s734_val_n3;
    end
    always @(posedge \clk ) begin
        s735_val_n4 <= s734_val_n4;
    end
    always @(posedge \clk ) begin
        s735_val_n5 <= s734_val_n5;
    end
    always @(posedge \clk ) begin
        s735_val_n6 <= s734_val_n6;
    end
    always @(posedge \clk ) begin
        s735_val_n7 <= s734_val_n7;
    end
    always @(posedge \clk ) begin
        \s736_val  <= \s735_val ;
    end
    always @(posedge \clk ) begin
        s736_val_n1 <= s735_val_n1;
    end
    always @(posedge \clk ) begin
        s736_val_n2 <= s735_val_n2;
    end
    always @(posedge \clk ) begin
        s736_val_n3 <= s735_val_n3;
    end
    always @(posedge \clk ) begin
        s736_val_n4 <= s735_val_n4;
    end
    always @(posedge \clk ) begin
        s736_val_n5 <= s735_val_n5;
    end
    always @(posedge \clk ) begin
        s736_val_n6 <= s735_val_n6;
    end
    always @(posedge \clk ) begin
        s736_val_n7 <= s735_val_n7;
    end
    always @(posedge \clk ) begin
        \s737_val  <= \s736_val ;
    end
    always @(posedge \clk ) begin
        s737_val_n1 <= s736_val_n1;
    end
    always @(posedge \clk ) begin
        s737_val_n2 <= s736_val_n2;
    end
    always @(posedge \clk ) begin
        s737_val_n3 <= s736_val_n3;
    end
    always @(posedge \clk ) begin
        s737_val_n4 <= s736_val_n4;
    end
    always @(posedge \clk ) begin
        s737_val_n5 <= s736_val_n5;
    end
    always @(posedge \clk ) begin
        s737_val_n6 <= s736_val_n6;
    end
    always @(posedge \clk ) begin
        s737_val_n7 <= s736_val_n7;
    end
    always @(posedge \clk ) begin
        \s738_val  <= \s737_val ;
    end
    always @(posedge \clk ) begin
        s738_val_n1 <= s737_val_n1;
    end
    always @(posedge \clk ) begin
        s738_val_n2 <= s737_val_n2;
    end
    always @(posedge \clk ) begin
        s738_val_n3 <= s737_val_n3;
    end
    always @(posedge \clk ) begin
        s738_val_n4 <= s737_val_n4;
    end
    always @(posedge \clk ) begin
        s738_val_n5 <= s737_val_n5;
    end
    always @(posedge \clk ) begin
        s738_val_n6 <= s737_val_n6;
    end
    always @(posedge \clk ) begin
        s738_val_n7 <= s737_val_n7;
    end
    always @(posedge \clk ) begin
        \s739_val  <= \s738_val ;
    end
    always @(posedge \clk ) begin
        s739_val_n1 <= s738_val_n1;
    end
    always @(posedge \clk ) begin
        s739_val_n2 <= s738_val_n2;
    end
    always @(posedge \clk ) begin
        s739_val_n3 <= s738_val_n3;
    end
    always @(posedge \clk ) begin
        s739_val_n4 <= s738_val_n4;
    end
    always @(posedge \clk ) begin
        s739_val_n5 <= s738_val_n5;
    end
    always @(posedge \clk ) begin
        s739_val_n6 <= s738_val_n6;
    end
    always @(posedge \clk ) begin
        s739_val_n7 <= s738_val_n7;
    end
    always @(posedge \clk ) begin
        \s740_val  <= \s739_val ;
    end
    always @(posedge \clk ) begin
        s740_val_n1 <= s739_val_n1;
    end
    always @(posedge \clk ) begin
        s740_val_n2 <= s739_val_n2;
    end
    always @(posedge \clk ) begin
        s740_val_n3 <= s739_val_n3;
    end
    always @(posedge \clk ) begin
        s740_val_n4 <= s739_val_n4;
    end
    always @(posedge \clk ) begin
        s740_val_n5 <= s739_val_n5;
    end
    always @(posedge \clk ) begin
        s740_val_n6 <= s739_val_n6;
    end
    always @(posedge \clk ) begin
        s740_val_n7 <= s739_val_n7;
    end
    always @(posedge \clk ) begin
        \s741_val  <= \s740_val ;
    end
    always @(posedge \clk ) begin
        s741_val_n1 <= s740_val_n1;
    end
    always @(posedge \clk ) begin
        s741_val_n2 <= s740_val_n2;
    end
    always @(posedge \clk ) begin
        s741_val_n3 <= s740_val_n3;
    end
    always @(posedge \clk ) begin
        s741_val_n4 <= s740_val_n4;
    end
    always @(posedge \clk ) begin
        s741_val_n5 <= s740_val_n5;
    end
    always @(posedge \clk ) begin
        s741_val_n6 <= s740_val_n6;
    end
    always @(posedge \clk ) begin
        s741_val_n7 <= s740_val_n7;
    end
    always @(posedge \clk ) begin
        \s742_val  <= \s741_val ;
    end
    always @(posedge \clk ) begin
        s742_val_n1 <= s741_val_n1;
    end
    always @(posedge \clk ) begin
        s742_val_n2 <= s741_val_n2;
    end
    always @(posedge \clk ) begin
        s742_val_n3 <= s741_val_n3;
    end
    always @(posedge \clk ) begin
        s742_val_n4 <= s741_val_n4;
    end
    always @(posedge \clk ) begin
        s742_val_n5 <= s741_val_n5;
    end
    always @(posedge \clk ) begin
        s742_val_n6 <= s741_val_n6;
    end
    always @(posedge \clk ) begin
        s742_val_n7 <= s741_val_n7;
    end
    always @(posedge \clk ) begin
        \s743_val  <= \s742_val ;
    end
    always @(posedge \clk ) begin
        s743_val_n1 <= s742_val_n1;
    end
    always @(posedge \clk ) begin
        s743_val_n2 <= s742_val_n2;
    end
    always @(posedge \clk ) begin
        s743_val_n3 <= s742_val_n3;
    end
    always @(posedge \clk ) begin
        s743_val_n4 <= s742_val_n4;
    end
    always @(posedge \clk ) begin
        s743_val_n5 <= s742_val_n5;
    end
    always @(posedge \clk ) begin
        s743_val_n6 <= s742_val_n6;
    end
    always @(posedge \clk ) begin
        s743_val_n7 <= s742_val_n7;
    end
    always @(posedge \clk ) begin
        \s744_val  <= \s743_val ;
    end
    always @(posedge \clk ) begin
        s744_val_n1 <= s743_val_n1;
    end
    always @(posedge \clk ) begin
        s744_val_n2 <= s743_val_n2;
    end
    always @(posedge \clk ) begin
        s744_val_n3 <= s743_val_n3;
    end
    always @(posedge \clk ) begin
        s744_val_n4 <= s743_val_n4;
    end
    always @(posedge \clk ) begin
        s744_val_n5 <= s743_val_n5;
    end
    always @(posedge \clk ) begin
        s744_val_n6 <= s743_val_n6;
    end
    always @(posedge \clk ) begin
        s744_val_n7 <= s743_val_n7;
    end
    always @(posedge \clk ) begin
        \s745_val  <= \s744_val ;
    end
    always @(posedge \clk ) begin
        s745_val_n1 <= s744_val_n1;
    end
    always @(posedge \clk ) begin
        s745_val_n2 <= s744_val_n2;
    end
    always @(posedge \clk ) begin
        s745_val_n3 <= s744_val_n3;
    end
    always @(posedge \clk ) begin
        s745_val_n4 <= s744_val_n4;
    end
    always @(posedge \clk ) begin
        s745_val_n5 <= s744_val_n5;
    end
    always @(posedge \clk ) begin
        s745_val_n6 <= s744_val_n6;
    end
    always @(posedge \clk ) begin
        s745_val_n7 <= s744_val_n7;
    end
    always @(posedge \clk ) begin
        \s746_val  <= \s745_val ;
    end
    always @(posedge \clk ) begin
        s746_val_n1 <= s745_val_n1;
    end
    always @(posedge \clk ) begin
        s746_val_n2 <= s745_val_n2;
    end
    always @(posedge \clk ) begin
        s746_val_n3 <= s745_val_n3;
    end
    always @(posedge \clk ) begin
        s746_val_n4 <= s745_val_n4;
    end
    always @(posedge \clk ) begin
        s746_val_n5 <= s745_val_n5;
    end
    always @(posedge \clk ) begin
        s746_val_n6 <= s745_val_n6;
    end
    always @(posedge \clk ) begin
        s746_val_n7 <= s745_val_n7;
    end
    always @(posedge \clk ) begin
        \s747_val  <= \s746_val ;
    end
    always @(posedge \clk ) begin
        s747_val_n1 <= s746_val_n1;
    end
    always @(posedge \clk ) begin
        s747_val_n2 <= s746_val_n2;
    end
    always @(posedge \clk ) begin
        s747_val_n3 <= s746_val_n3;
    end
    always @(posedge \clk ) begin
        s747_val_n4 <= s746_val_n4;
    end
    always @(posedge \clk ) begin
        s747_val_n5 <= s746_val_n5;
    end
    always @(posedge \clk ) begin
        s747_val_n6 <= s746_val_n6;
    end
    always @(posedge \clk ) begin
        s747_val_n7 <= s746_val_n7;
    end
    always @(posedge \clk ) begin
        \s748_val  <= \s747_val ;
    end
    always @(posedge \clk ) begin
        s748_val_n1 <= s747_val_n1;
    end
    always @(posedge \clk ) begin
        s748_val_n2 <= s747_val_n2;
    end
    always @(posedge \clk ) begin
        s748_val_n3 <= s747_val_n3;
    end
    always @(posedge \clk ) begin
        s748_val_n4 <= s747_val_n4;
    end
    always @(posedge \clk ) begin
        s748_val_n5 <= s747_val_n5;
    end
    always @(posedge \clk ) begin
        s748_val_n6 <= s747_val_n6;
    end
    always @(posedge \clk ) begin
        s748_val_n7 <= s747_val_n7;
    end
    always @(posedge \clk ) begin
        \s749_val  <= \s748_val ;
    end
    always @(posedge \clk ) begin
        s749_val_n1 <= s748_val_n1;
    end
    always @(posedge \clk ) begin
        s749_val_n2 <= s748_val_n2;
    end
    always @(posedge \clk ) begin
        s749_val_n3 <= s748_val_n3;
    end
    always @(posedge \clk ) begin
        s749_val_n4 <= s748_val_n4;
    end
    always @(posedge \clk ) begin
        s749_val_n5 <= s748_val_n5;
    end
    always @(posedge \clk ) begin
        s749_val_n6 <= s748_val_n6;
    end
    always @(posedge \clk ) begin
        s749_val_n7 <= s748_val_n7;
    end
    always @(posedge \clk ) begin
        \s750_val  <= \s749_val ;
    end
    always @(posedge \clk ) begin
        s750_val_n1 <= s749_val_n1;
    end
    always @(posedge \clk ) begin
        s750_val_n2 <= s749_val_n2;
    end
    always @(posedge \clk ) begin
        s750_val_n3 <= s749_val_n3;
    end
    always @(posedge \clk ) begin
        s750_val_n4 <= s749_val_n4;
    end
    always @(posedge \clk ) begin
        s750_val_n5 <= s749_val_n5;
    end
    always @(posedge \clk ) begin
        s750_val_n6 <= s749_val_n6;
    end
    always @(posedge \clk ) begin
        s750_val_n7 <= s749_val_n7;
    end
    always @(posedge \clk ) begin
        \s751_val  <= \s750_val ;
    end
    always @(posedge \clk ) begin
        s751_val_n1 <= s750_val_n1;
    end
    always @(posedge \clk ) begin
        s751_val_n2 <= s750_val_n2;
    end
    always @(posedge \clk ) begin
        s751_val_n3 <= s750_val_n3;
    end
    always @(posedge \clk ) begin
        s751_val_n4 <= s750_val_n4;
    end
    always @(posedge \clk ) begin
        s751_val_n5 <= s750_val_n5;
    end
    always @(posedge \clk ) begin
        s751_val_n6 <= s750_val_n6;
    end
    always @(posedge \clk ) begin
        s751_val_n7 <= s750_val_n7;
    end
    always @(posedge \clk ) begin
        \s752_val  <= \s751_val ;
    end
    always @(posedge \clk ) begin
        s752_val_n1 <= s751_val_n1;
    end
    always @(posedge \clk ) begin
        s752_val_n2 <= s751_val_n2;
    end
    always @(posedge \clk ) begin
        s752_val_n3 <= s751_val_n3;
    end
    always @(posedge \clk ) begin
        s752_val_n4 <= s751_val_n4;
    end
    always @(posedge \clk ) begin
        s752_val_n5 <= s751_val_n5;
    end
    always @(posedge \clk ) begin
        s752_val_n6 <= s751_val_n6;
    end
    always @(posedge \clk ) begin
        s752_val_n7 <= s751_val_n7;
    end
    always @(posedge \clk ) begin
        \s753_val  <= \s752_val ;
    end
    always @(posedge \clk ) begin
        s753_val_n1 <= s752_val_n1;
    end
    always @(posedge \clk ) begin
        s753_val_n2 <= s752_val_n2;
    end
    always @(posedge \clk ) begin
        s753_val_n3 <= s752_val_n3;
    end
    always @(posedge \clk ) begin
        s753_val_n4 <= s752_val_n4;
    end
    always @(posedge \clk ) begin
        s753_val_n5 <= s752_val_n5;
    end
    always @(posedge \clk ) begin
        s753_val_n6 <= s752_val_n6;
    end
    always @(posedge \clk ) begin
        s753_val_n7 <= s752_val_n7;
    end
    always @(posedge \clk ) begin
        \s754_val  <= \s753_val ;
    end
    always @(posedge \clk ) begin
        s754_val_n1 <= s753_val_n1;
    end
    always @(posedge \clk ) begin
        s754_val_n2 <= s753_val_n2;
    end
    always @(posedge \clk ) begin
        s754_val_n3 <= s753_val_n3;
    end
    always @(posedge \clk ) begin
        s754_val_n4 <= s753_val_n4;
    end
    always @(posedge \clk ) begin
        s754_val_n5 <= s753_val_n5;
    end
    always @(posedge \clk ) begin
        s754_val_n6 <= s753_val_n6;
    end
    always @(posedge \clk ) begin
        s754_val_n7 <= s753_val_n7;
    end
    always @(posedge \clk ) begin
        \s755_val  <= \s754_val ;
    end
    always @(posedge \clk ) begin
        s755_val_n1 <= s754_val_n1;
    end
    always @(posedge \clk ) begin
        s755_val_n2 <= s754_val_n2;
    end
    always @(posedge \clk ) begin
        s755_val_n3 <= s754_val_n3;
    end
    always @(posedge \clk ) begin
        s755_val_n4 <= s754_val_n4;
    end
    always @(posedge \clk ) begin
        s755_val_n5 <= s754_val_n5;
    end
    always @(posedge \clk ) begin
        s755_val_n6 <= s754_val_n6;
    end
    always @(posedge \clk ) begin
        s755_val_n7 <= s754_val_n7;
    end
    always @(posedge \clk ) begin
        \s756_val  <= \s755_val ;
    end
    always @(posedge \clk ) begin
        s756_val_n1 <= s755_val_n1;
    end
    always @(posedge \clk ) begin
        s756_val_n2 <= s755_val_n2;
    end
    always @(posedge \clk ) begin
        s756_val_n3 <= s755_val_n3;
    end
    always @(posedge \clk ) begin
        s756_val_n4 <= s755_val_n4;
    end
    always @(posedge \clk ) begin
        s756_val_n5 <= s755_val_n5;
    end
    always @(posedge \clk ) begin
        s756_val_n6 <= s755_val_n6;
    end
    always @(posedge \clk ) begin
        s756_val_n7 <= s755_val_n7;
    end
    always @(posedge \clk ) begin
        \s757_val  <= \s756_val ;
    end
    always @(posedge \clk ) begin
        s757_val_n1 <= s756_val_n1;
    end
    always @(posedge \clk ) begin
        s757_val_n2 <= s756_val_n2;
    end
    always @(posedge \clk ) begin
        s757_val_n3 <= s756_val_n3;
    end
    always @(posedge \clk ) begin
        s757_val_n4 <= s756_val_n4;
    end
    always @(posedge \clk ) begin
        s757_val_n5 <= s756_val_n5;
    end
    always @(posedge \clk ) begin
        s757_val_n6 <= s756_val_n6;
    end
    always @(posedge \clk ) begin
        s757_val_n7 <= s756_val_n7;
    end
    always @(posedge \clk ) begin
        \s758_val  <= \s757_val ;
    end
    always @(posedge \clk ) begin
        s758_val_n1 <= s757_val_n1;
    end
    always @(posedge \clk ) begin
        s758_val_n2 <= s757_val_n2;
    end
    always @(posedge \clk ) begin
        s758_val_n3 <= s757_val_n3;
    end
    always @(posedge \clk ) begin
        s758_val_n4 <= s757_val_n4;
    end
    always @(posedge \clk ) begin
        s758_val_n5 <= s757_val_n5;
    end
    always @(posedge \clk ) begin
        s758_val_n6 <= s757_val_n6;
    end
    always @(posedge \clk ) begin
        s758_val_n7 <= s757_val_n7;
    end
    always @(posedge \clk ) begin
        \s759_val  <= \s758_val ;
    end
    always @(posedge \clk ) begin
        s759_val_n1 <= s758_val_n1;
    end
    always @(posedge \clk ) begin
        s759_val_n2 <= s758_val_n2;
    end
    always @(posedge \clk ) begin
        s759_val_n3 <= s758_val_n3;
    end
    always @(posedge \clk ) begin
        s759_val_n4 <= s758_val_n4;
    end
    always @(posedge \clk ) begin
        s759_val_n5 <= s758_val_n5;
    end
    always @(posedge \clk ) begin
        s759_val_n6 <= s758_val_n6;
    end
    always @(posedge \clk ) begin
        s759_val_n7 <= s758_val_n7;
    end
    always @(posedge \clk ) begin
        \s760_val  <= \s759_val ;
    end
    always @(posedge \clk ) begin
        s760_val_n1 <= s759_val_n1;
    end
    always @(posedge \clk ) begin
        s760_val_n2 <= s759_val_n2;
    end
    always @(posedge \clk ) begin
        s760_val_n3 <= s759_val_n3;
    end
    always @(posedge \clk ) begin
        s760_val_n4 <= s759_val_n4;
    end
    always @(posedge \clk ) begin
        s760_val_n5 <= s759_val_n5;
    end
    always @(posedge \clk ) begin
        s760_val_n6 <= s759_val_n6;
    end
    always @(posedge \clk ) begin
        s760_val_n7 <= s759_val_n7;
    end
    always @(posedge \clk ) begin
        \s761_val  <= \s760_val ;
    end
    always @(posedge \clk ) begin
        s761_val_n1 <= s760_val_n1;
    end
    always @(posedge \clk ) begin
        s761_val_n2 <= s760_val_n2;
    end
    always @(posedge \clk ) begin
        s761_val_n3 <= s760_val_n3;
    end
    always @(posedge \clk ) begin
        s761_val_n4 <= s760_val_n4;
    end
    always @(posedge \clk ) begin
        s761_val_n5 <= s760_val_n5;
    end
    always @(posedge \clk ) begin
        s761_val_n6 <= s760_val_n6;
    end
    always @(posedge \clk ) begin
        s761_val_n7 <= s760_val_n7;
    end
    always @(posedge \clk ) begin
        \s762_val  <= \s761_val ;
    end
    always @(posedge \clk ) begin
        s762_val_n1 <= s761_val_n1;
    end
    always @(posedge \clk ) begin
        s762_val_n2 <= s761_val_n2;
    end
    always @(posedge \clk ) begin
        s762_val_n3 <= s761_val_n3;
    end
    always @(posedge \clk ) begin
        s762_val_n4 <= s761_val_n4;
    end
    always @(posedge \clk ) begin
        s762_val_n5 <= s761_val_n5;
    end
    always @(posedge \clk ) begin
        s762_val_n6 <= s761_val_n6;
    end
    always @(posedge \clk ) begin
        s762_val_n7 <= s761_val_n7;
    end
    always @(posedge \clk ) begin
        \s763_val  <= \s762_val ;
    end
    always @(posedge \clk ) begin
        s763_val_n1 <= s762_val_n1;
    end
    always @(posedge \clk ) begin
        s763_val_n2 <= s762_val_n2;
    end
    always @(posedge \clk ) begin
        s763_val_n3 <= s762_val_n3;
    end
    always @(posedge \clk ) begin
        s763_val_n4 <= s762_val_n4;
    end
    always @(posedge \clk ) begin
        s763_val_n5 <= s762_val_n5;
    end
    always @(posedge \clk ) begin
        s763_val_n6 <= s762_val_n6;
    end
    always @(posedge \clk ) begin
        s763_val_n7 <= s762_val_n7;
    end
    always @(posedge \clk ) begin
        \s764_val  <= \s763_val ;
    end
    always @(posedge \clk ) begin
        s764_val_n1 <= s763_val_n1;
    end
    always @(posedge \clk ) begin
        s764_val_n2 <= s763_val_n2;
    end
    always @(posedge \clk ) begin
        s764_val_n3 <= s763_val_n3;
    end
    always @(posedge \clk ) begin
        s764_val_n4 <= s763_val_n4;
    end
    always @(posedge \clk ) begin
        s764_val_n5 <= s763_val_n5;
    end
    always @(posedge \clk ) begin
        s764_val_n6 <= s763_val_n6;
    end
    always @(posedge \clk ) begin
        s764_val_n7 <= s763_val_n7;
    end
    always @(posedge \clk ) begin
        \s765_val  <= \s764_val ;
    end
    always @(posedge \clk ) begin
        s765_val_n1 <= s764_val_n1;
    end
    always @(posedge \clk ) begin
        s765_val_n2 <= s764_val_n2;
    end
    always @(posedge \clk ) begin
        s765_val_n3 <= s764_val_n3;
    end
    always @(posedge \clk ) begin
        s765_val_n4 <= s764_val_n4;
    end
    always @(posedge \clk ) begin
        s765_val_n5 <= s764_val_n5;
    end
    always @(posedge \clk ) begin
        s765_val_n6 <= s764_val_n6;
    end
    always @(posedge \clk ) begin
        s765_val_n7 <= s764_val_n7;
    end
    always @(posedge \clk ) begin
        \s766_val  <= \s765_val ;
    end
    always @(posedge \clk ) begin
        s766_val_n1 <= s765_val_n1;
    end
    always @(posedge \clk ) begin
        s766_val_n2 <= s765_val_n2;
    end
    always @(posedge \clk ) begin
        s766_val_n3 <= s765_val_n3;
    end
    always @(posedge \clk ) begin
        s766_val_n4 <= s765_val_n4;
    end
    always @(posedge \clk ) begin
        s766_val_n5 <= s765_val_n5;
    end
    always @(posedge \clk ) begin
        s766_val_n6 <= s765_val_n6;
    end
    always @(posedge \clk ) begin
        s766_val_n7 <= s765_val_n7;
    end
    always @(posedge \clk ) begin
        \s767_val  <= \s766_val ;
    end
    always @(posedge \clk ) begin
        s767_val_n1 <= s766_val_n1;
    end
    always @(posedge \clk ) begin
        s767_val_n2 <= s766_val_n2;
    end
    always @(posedge \clk ) begin
        s767_val_n3 <= s766_val_n3;
    end
    always @(posedge \clk ) begin
        s767_val_n4 <= s766_val_n4;
    end
    always @(posedge \clk ) begin
        s767_val_n5 <= s766_val_n5;
    end
    always @(posedge \clk ) begin
        s767_val_n6 <= s766_val_n6;
    end
    always @(posedge \clk ) begin
        s767_val_n7 <= s766_val_n7;
    end
    always @(posedge \clk ) begin
        \s768_val  <= \s767_val ;
    end
    always @(posedge \clk ) begin
        s768_val_n1 <= s767_val_n1;
    end
    always @(posedge \clk ) begin
        s768_val_n2 <= s767_val_n2;
    end
    always @(posedge \clk ) begin
        s768_val_n3 <= s767_val_n3;
    end
    always @(posedge \clk ) begin
        s768_val_n4 <= s767_val_n4;
    end
    always @(posedge \clk ) begin
        s768_val_n5 <= s767_val_n5;
    end
    always @(posedge \clk ) begin
        s768_val_n6 <= s767_val_n6;
    end
    always @(posedge \clk ) begin
        s768_val_n7 <= s767_val_n7;
    end
    always @(posedge \clk ) begin
        \s769_val  <= \s768_val ;
    end
    always @(posedge \clk ) begin
        s769_val_n1 <= s768_val_n1;
    end
    always @(posedge \clk ) begin
        s769_val_n2 <= s768_val_n2;
    end
    always @(posedge \clk ) begin
        s769_val_n3 <= s768_val_n3;
    end
    always @(posedge \clk ) begin
        s769_val_n4 <= s768_val_n4;
    end
    always @(posedge \clk ) begin
        s769_val_n5 <= s768_val_n5;
    end
    always @(posedge \clk ) begin
        s769_val_n6 <= s768_val_n6;
    end
    always @(posedge \clk ) begin
        s769_val_n7 <= s768_val_n7;
    end
    always @(posedge \clk ) begin
        \s770_val  <= \s769_val ;
    end
    always @(posedge \clk ) begin
        s770_val_n1 <= s769_val_n1;
    end
    always @(posedge \clk ) begin
        s770_val_n2 <= s769_val_n2;
    end
    always @(posedge \clk ) begin
        s770_val_n3 <= s769_val_n3;
    end
    always @(posedge \clk ) begin
        s770_val_n4 <= s769_val_n4;
    end
    always @(posedge \clk ) begin
        s770_val_n5 <= s769_val_n5;
    end
    always @(posedge \clk ) begin
        s770_val_n6 <= s769_val_n6;
    end
    always @(posedge \clk ) begin
        s770_val_n7 <= s769_val_n7;
    end
    always @(posedge \clk ) begin
        \s771_val  <= \s770_val ;
    end
    always @(posedge \clk ) begin
        s771_val_n1 <= s770_val_n1;
    end
    always @(posedge \clk ) begin
        s771_val_n2 <= s770_val_n2;
    end
    always @(posedge \clk ) begin
        s771_val_n3 <= s770_val_n3;
    end
    always @(posedge \clk ) begin
        s771_val_n4 <= s770_val_n4;
    end
    always @(posedge \clk ) begin
        s771_val_n5 <= s770_val_n5;
    end
    always @(posedge \clk ) begin
        s771_val_n6 <= s770_val_n6;
    end
    always @(posedge \clk ) begin
        s771_val_n7 <= s770_val_n7;
    end
    always @(posedge \clk ) begin
        \s772_val  <= \s771_val ;
    end
    always @(posedge \clk ) begin
        s772_val_n1 <= s771_val_n1;
    end
    always @(posedge \clk ) begin
        s772_val_n2 <= s771_val_n2;
    end
    always @(posedge \clk ) begin
        s772_val_n3 <= s771_val_n3;
    end
    always @(posedge \clk ) begin
        s772_val_n4 <= s771_val_n4;
    end
    always @(posedge \clk ) begin
        s772_val_n5 <= s771_val_n5;
    end
    always @(posedge \clk ) begin
        s772_val_n6 <= s771_val_n6;
    end
    always @(posedge \clk ) begin
        s772_val_n7 <= s771_val_n7;
    end
    always @(posedge \clk ) begin
        \s773_val  <= \s772_val ;
    end
    always @(posedge \clk ) begin
        s773_val_n1 <= s772_val_n1;
    end
    always @(posedge \clk ) begin
        s773_val_n2 <= s772_val_n2;
    end
    always @(posedge \clk ) begin
        s773_val_n3 <= s772_val_n3;
    end
    always @(posedge \clk ) begin
        s773_val_n4 <= s772_val_n4;
    end
    always @(posedge \clk ) begin
        s773_val_n5 <= s772_val_n5;
    end
    always @(posedge \clk ) begin
        s773_val_n6 <= s772_val_n6;
    end
    always @(posedge \clk ) begin
        s773_val_n7 <= s772_val_n7;
    end
    always @(posedge \clk ) begin
        \s774_val  <= \s773_val ;
    end
    always @(posedge \clk ) begin
        s774_val_n1 <= s773_val_n1;
    end
    always @(posedge \clk ) begin
        s774_val_n2 <= s773_val_n2;
    end
    always @(posedge \clk ) begin
        s774_val_n3 <= s773_val_n3;
    end
    always @(posedge \clk ) begin
        s774_val_n4 <= s773_val_n4;
    end
    always @(posedge \clk ) begin
        s774_val_n5 <= s773_val_n5;
    end
    always @(posedge \clk ) begin
        s774_val_n6 <= s773_val_n6;
    end
    always @(posedge \clk ) begin
        s774_val_n7 <= s773_val_n7;
    end
    always @(posedge \clk ) begin
        \s775_val  <= \s774_val ;
    end
    always @(posedge \clk ) begin
        s775_val_n1 <= s774_val_n1;
    end
    always @(posedge \clk ) begin
        s775_val_n2 <= s774_val_n2;
    end
    always @(posedge \clk ) begin
        s775_val_n3 <= s774_val_n3;
    end
    always @(posedge \clk ) begin
        s775_val_n4 <= s774_val_n4;
    end
    always @(posedge \clk ) begin
        s775_val_n5 <= s774_val_n5;
    end
    always @(posedge \clk ) begin
        s775_val_n6 <= s774_val_n6;
    end
    always @(posedge \clk ) begin
        s775_val_n7 <= s774_val_n7;
    end
    always @(posedge \clk ) begin
        \s776_val  <= \s775_val ;
    end
    always @(posedge \clk ) begin
        s776_val_n1 <= s775_val_n1;
    end
    always @(posedge \clk ) begin
        s776_val_n2 <= s775_val_n2;
    end
    always @(posedge \clk ) begin
        s776_val_n3 <= s775_val_n3;
    end
    always @(posedge \clk ) begin
        s776_val_n4 <= s775_val_n4;
    end
    always @(posedge \clk ) begin
        s776_val_n5 <= s775_val_n5;
    end
    always @(posedge \clk ) begin
        s776_val_n6 <= s775_val_n6;
    end
    always @(posedge \clk ) begin
        s776_val_n7 <= s775_val_n7;
    end
    always @(posedge \clk ) begin
        \s777_val  <= \s776_val ;
    end
    always @(posedge \clk ) begin
        s777_val_n1 <= s776_val_n1;
    end
    always @(posedge \clk ) begin
        s777_val_n2 <= s776_val_n2;
    end
    always @(posedge \clk ) begin
        s777_val_n3 <= s776_val_n3;
    end
    always @(posedge \clk ) begin
        s777_val_n4 <= s776_val_n4;
    end
    always @(posedge \clk ) begin
        s777_val_n5 <= s776_val_n5;
    end
    always @(posedge \clk ) begin
        s777_val_n6 <= s776_val_n6;
    end
    always @(posedge \clk ) begin
        s777_val_n7 <= s776_val_n7;
    end
    always @(posedge \clk ) begin
        \s778_val  <= \s777_val ;
    end
    always @(posedge \clk ) begin
        s778_val_n1 <= s777_val_n1;
    end
    always @(posedge \clk ) begin
        s778_val_n2 <= s777_val_n2;
    end
    always @(posedge \clk ) begin
        s778_val_n3 <= s777_val_n3;
    end
    always @(posedge \clk ) begin
        s778_val_n4 <= s777_val_n4;
    end
    always @(posedge \clk ) begin
        s778_val_n5 <= s777_val_n5;
    end
    always @(posedge \clk ) begin
        s778_val_n6 <= s777_val_n6;
    end
    always @(posedge \clk ) begin
        s778_val_n7 <= s777_val_n7;
    end
    always @(posedge \clk ) begin
        \s779_val  <= \s778_val ;
    end
    always @(posedge \clk ) begin
        s779_val_n1 <= s778_val_n1;
    end
    always @(posedge \clk ) begin
        s779_val_n2 <= s778_val_n2;
    end
    always @(posedge \clk ) begin
        s779_val_n3 <= s778_val_n3;
    end
    always @(posedge \clk ) begin
        s779_val_n4 <= s778_val_n4;
    end
    always @(posedge \clk ) begin
        s779_val_n5 <= s778_val_n5;
    end
    always @(posedge \clk ) begin
        s779_val_n6 <= s778_val_n6;
    end
    always @(posedge \clk ) begin
        s779_val_n7 <= s778_val_n7;
    end
    always @(posedge \clk ) begin
        \s780_val  <= \s779_val ;
    end
    always @(posedge \clk ) begin
        s780_val_n1 <= s779_val_n1;
    end
    always @(posedge \clk ) begin
        s780_val_n2 <= s779_val_n2;
    end
    always @(posedge \clk ) begin
        s780_val_n3 <= s779_val_n3;
    end
    always @(posedge \clk ) begin
        s780_val_n4 <= s779_val_n4;
    end
    always @(posedge \clk ) begin
        s780_val_n5 <= s779_val_n5;
    end
    always @(posedge \clk ) begin
        s780_val_n6 <= s779_val_n6;
    end
    always @(posedge \clk ) begin
        s780_val_n7 <= s779_val_n7;
    end
    always @(posedge \clk ) begin
        \s781_val  <= \s780_val ;
    end
    always @(posedge \clk ) begin
        s781_val_n1 <= s780_val_n1;
    end
    always @(posedge \clk ) begin
        s781_val_n2 <= s780_val_n2;
    end
    always @(posedge \clk ) begin
        s781_val_n3 <= s780_val_n3;
    end
    always @(posedge \clk ) begin
        s781_val_n4 <= s780_val_n4;
    end
    always @(posedge \clk ) begin
        s781_val_n5 <= s780_val_n5;
    end
    always @(posedge \clk ) begin
        s781_val_n6 <= s780_val_n6;
    end
    always @(posedge \clk ) begin
        s781_val_n7 <= s780_val_n7;
    end
    always @(posedge \clk ) begin
        \s782_val  <= \s781_val ;
    end
    always @(posedge \clk ) begin
        s782_val_n1 <= s781_val_n1;
    end
    always @(posedge \clk ) begin
        s782_val_n2 <= s781_val_n2;
    end
    always @(posedge \clk ) begin
        s782_val_n3 <= s781_val_n3;
    end
    always @(posedge \clk ) begin
        s782_val_n4 <= s781_val_n4;
    end
    always @(posedge \clk ) begin
        s782_val_n5 <= s781_val_n5;
    end
    always @(posedge \clk ) begin
        s782_val_n6 <= s781_val_n6;
    end
    always @(posedge \clk ) begin
        s782_val_n7 <= s781_val_n7;
    end
    always @(posedge \clk ) begin
        \s783_val  <= \s782_val ;
    end
    always @(posedge \clk ) begin
        s783_val_n1 <= s782_val_n1;
    end
    always @(posedge \clk ) begin
        s783_val_n2 <= s782_val_n2;
    end
    always @(posedge \clk ) begin
        s783_val_n3 <= s782_val_n3;
    end
    always @(posedge \clk ) begin
        s783_val_n4 <= s782_val_n4;
    end
    always @(posedge \clk ) begin
        s783_val_n5 <= s782_val_n5;
    end
    always @(posedge \clk ) begin
        s783_val_n6 <= s782_val_n6;
    end
    always @(posedge \clk ) begin
        s783_val_n7 <= s782_val_n7;
    end
    always @(posedge \clk ) begin
        \s784_val  <= \s783_val ;
    end
    always @(posedge \clk ) begin
        s784_val_n1 <= s783_val_n1;
    end
    always @(posedge \clk ) begin
        s784_val_n2 <= s783_val_n2;
    end
    always @(posedge \clk ) begin
        s784_val_n3 <= s783_val_n3;
    end
    always @(posedge \clk ) begin
        s784_val_n4 <= s783_val_n4;
    end
    always @(posedge \clk ) begin
        s784_val_n5 <= s783_val_n5;
    end
    always @(posedge \clk ) begin
        s784_val_n6 <= s783_val_n6;
    end
    always @(posedge \clk ) begin
        s784_val_n7 <= s783_val_n7;
    end
    always @(posedge \clk ) begin
        \s785_val  <= \s784_val ;
    end
    always @(posedge \clk ) begin
        s785_val_n1 <= s784_val_n1;
    end
    always @(posedge \clk ) begin
        s785_val_n2 <= s784_val_n2;
    end
    always @(posedge \clk ) begin
        s785_val_n3 <= s784_val_n3;
    end
    always @(posedge \clk ) begin
        s785_val_n4 <= s784_val_n4;
    end
    always @(posedge \clk ) begin
        s785_val_n5 <= s784_val_n5;
    end
    always @(posedge \clk ) begin
        s785_val_n6 <= s784_val_n6;
    end
    always @(posedge \clk ) begin
        s785_val_n7 <= s784_val_n7;
    end
    always @(posedge \clk ) begin
        \s786_val  <= \s785_val ;
    end
    always @(posedge \clk ) begin
        s786_val_n1 <= s785_val_n1;
    end
    always @(posedge \clk ) begin
        s786_val_n2 <= s785_val_n2;
    end
    always @(posedge \clk ) begin
        s786_val_n3 <= s785_val_n3;
    end
    always @(posedge \clk ) begin
        s786_val_n4 <= s785_val_n4;
    end
    always @(posedge \clk ) begin
        s786_val_n5 <= s785_val_n5;
    end
    always @(posedge \clk ) begin
        s786_val_n6 <= s785_val_n6;
    end
    always @(posedge \clk ) begin
        s786_val_n7 <= s785_val_n7;
    end
    always @(posedge \clk ) begin
        \s787_val  <= \s786_val ;
    end
    always @(posedge \clk ) begin
        s787_val_n1 <= s786_val_n1;
    end
    always @(posedge \clk ) begin
        s787_val_n2 <= s786_val_n2;
    end
    always @(posedge \clk ) begin
        s787_val_n3 <= s786_val_n3;
    end
    always @(posedge \clk ) begin
        s787_val_n4 <= s786_val_n4;
    end
    always @(posedge \clk ) begin
        s787_val_n5 <= s786_val_n5;
    end
    always @(posedge \clk ) begin
        s787_val_n6 <= s786_val_n6;
    end
    always @(posedge \clk ) begin
        s787_val_n7 <= s786_val_n7;
    end
    always @(posedge \clk ) begin
        \s788_val  <= \s787_val ;
    end
    always @(posedge \clk ) begin
        s788_val_n1 <= s787_val_n1;
    end
    always @(posedge \clk ) begin
        s788_val_n2 <= s787_val_n2;
    end
    always @(posedge \clk ) begin
        s788_val_n3 <= s787_val_n3;
    end
    always @(posedge \clk ) begin
        s788_val_n4 <= s787_val_n4;
    end
    always @(posedge \clk ) begin
        s788_val_n5 <= s787_val_n5;
    end
    always @(posedge \clk ) begin
        s788_val_n6 <= s787_val_n6;
    end
    always @(posedge \clk ) begin
        s788_val_n7 <= s787_val_n7;
    end
    always @(posedge \clk ) begin
        \s789_val  <= \s788_val ;
    end
    always @(posedge \clk ) begin
        s789_val_n1 <= s788_val_n1;
    end
    always @(posedge \clk ) begin
        s789_val_n2 <= s788_val_n2;
    end
    always @(posedge \clk ) begin
        s789_val_n3 <= s788_val_n3;
    end
    always @(posedge \clk ) begin
        s789_val_n4 <= s788_val_n4;
    end
    always @(posedge \clk ) begin
        s789_val_n5 <= s788_val_n5;
    end
    always @(posedge \clk ) begin
        s789_val_n6 <= s788_val_n6;
    end
    always @(posedge \clk ) begin
        s789_val_n7 <= s788_val_n7;
    end
    always @(posedge \clk ) begin
        \s790_val  <= \s789_val ;
    end
    always @(posedge \clk ) begin
        s790_val_n1 <= s789_val_n1;
    end
    always @(posedge \clk ) begin
        s790_val_n2 <= s789_val_n2;
    end
    always @(posedge \clk ) begin
        s790_val_n3 <= s789_val_n3;
    end
    always @(posedge \clk ) begin
        s790_val_n4 <= s789_val_n4;
    end
    always @(posedge \clk ) begin
        s790_val_n5 <= s789_val_n5;
    end
    always @(posedge \clk ) begin
        s790_val_n6 <= s789_val_n6;
    end
    always @(posedge \clk ) begin
        s790_val_n7 <= s789_val_n7;
    end
    always @(posedge \clk ) begin
        \s791_val  <= \s790_val ;
    end
    always @(posedge \clk ) begin
        s791_val_n1 <= s790_val_n1;
    end
    always @(posedge \clk ) begin
        s791_val_n2 <= s790_val_n2;
    end
    always @(posedge \clk ) begin
        s791_val_n3 <= s790_val_n3;
    end
    always @(posedge \clk ) begin
        s791_val_n4 <= s790_val_n4;
    end
    always @(posedge \clk ) begin
        s791_val_n5 <= s790_val_n5;
    end
    always @(posedge \clk ) begin
        s791_val_n6 <= s790_val_n6;
    end
    always @(posedge \clk ) begin
        s791_val_n7 <= s790_val_n7;
    end
    always @(posedge \clk ) begin
        \s792_val  <= \s791_val ;
    end
    always @(posedge \clk ) begin
        s792_val_n1 <= s791_val_n1;
    end
    always @(posedge \clk ) begin
        s792_val_n2 <= s791_val_n2;
    end
    always @(posedge \clk ) begin
        s792_val_n3 <= s791_val_n3;
    end
    always @(posedge \clk ) begin
        s792_val_n4 <= s791_val_n4;
    end
    always @(posedge \clk ) begin
        s792_val_n5 <= s791_val_n5;
    end
    always @(posedge \clk ) begin
        s792_val_n6 <= s791_val_n6;
    end
    always @(posedge \clk ) begin
        s792_val_n7 <= s791_val_n7;
    end
    always @(posedge \clk ) begin
        \s793_val  <= \s792_val ;
    end
    always @(posedge \clk ) begin
        s793_val_n1 <= s792_val_n1;
    end
    always @(posedge \clk ) begin
        s793_val_n2 <= s792_val_n2;
    end
    always @(posedge \clk ) begin
        s793_val_n3 <= s792_val_n3;
    end
    always @(posedge \clk ) begin
        s793_val_n4 <= s792_val_n4;
    end
    always @(posedge \clk ) begin
        s793_val_n5 <= s792_val_n5;
    end
    always @(posedge \clk ) begin
        s793_val_n6 <= s792_val_n6;
    end
    always @(posedge \clk ) begin
        s793_val_n7 <= s792_val_n7;
    end
    always @(posedge \clk ) begin
        \s794_val  <= \s793_val ;
    end
    always @(posedge \clk ) begin
        s794_val_n1 <= s793_val_n1;
    end
    always @(posedge \clk ) begin
        s794_val_n2 <= s793_val_n2;
    end
    always @(posedge \clk ) begin
        s794_val_n3 <= s793_val_n3;
    end
    always @(posedge \clk ) begin
        s794_val_n4 <= s793_val_n4;
    end
    always @(posedge \clk ) begin
        s794_val_n5 <= s793_val_n5;
    end
    always @(posedge \clk ) begin
        s794_val_n6 <= s793_val_n6;
    end
    always @(posedge \clk ) begin
        s794_val_n7 <= s793_val_n7;
    end
    always @(posedge \clk ) begin
        \s795_val  <= \s794_val ;
    end
    always @(posedge \clk ) begin
        s795_val_n1 <= s794_val_n1;
    end
    always @(posedge \clk ) begin
        s795_val_n2 <= s794_val_n2;
    end
    always @(posedge \clk ) begin
        s795_val_n3 <= s794_val_n3;
    end
    always @(posedge \clk ) begin
        s795_val_n4 <= s794_val_n4;
    end
    always @(posedge \clk ) begin
        s795_val_n5 <= s794_val_n5;
    end
    always @(posedge \clk ) begin
        s795_val_n6 <= s794_val_n6;
    end
    always @(posedge \clk ) begin
        s795_val_n7 <= s794_val_n7;
    end
    always @(posedge \clk ) begin
        \s796_val  <= \s795_val ;
    end
    always @(posedge \clk ) begin
        s796_val_n1 <= s795_val_n1;
    end
    always @(posedge \clk ) begin
        s796_val_n2 <= s795_val_n2;
    end
    always @(posedge \clk ) begin
        s796_val_n3 <= s795_val_n3;
    end
    always @(posedge \clk ) begin
        s796_val_n4 <= s795_val_n4;
    end
    always @(posedge \clk ) begin
        s796_val_n5 <= s795_val_n5;
    end
    always @(posedge \clk ) begin
        s796_val_n6 <= s795_val_n6;
    end
    always @(posedge \clk ) begin
        s796_val_n7 <= s795_val_n7;
    end
    always @(posedge \clk ) begin
        \s797_val  <= \s796_val ;
    end
    always @(posedge \clk ) begin
        s797_val_n1 <= s796_val_n1;
    end
    always @(posedge \clk ) begin
        s797_val_n2 <= s796_val_n2;
    end
    always @(posedge \clk ) begin
        s797_val_n3 <= s796_val_n3;
    end
    always @(posedge \clk ) begin
        s797_val_n4 <= s796_val_n4;
    end
    always @(posedge \clk ) begin
        s797_val_n5 <= s796_val_n5;
    end
    always @(posedge \clk ) begin
        s797_val_n6 <= s796_val_n6;
    end
    always @(posedge \clk ) begin
        s797_val_n7 <= s796_val_n7;
    end
    always @(posedge \clk ) begin
        \s798_val  <= \s797_val ;
    end
    always @(posedge \clk ) begin
        s798_val_n1 <= s797_val_n1;
    end
    always @(posedge \clk ) begin
        s798_val_n2 <= s797_val_n2;
    end
    always @(posedge \clk ) begin
        s798_val_n3 <= s797_val_n3;
    end
    always @(posedge \clk ) begin
        s798_val_n4 <= s797_val_n4;
    end
    always @(posedge \clk ) begin
        s798_val_n5 <= s797_val_n5;
    end
    always @(posedge \clk ) begin
        s798_val_n6 <= s797_val_n6;
    end
    always @(posedge \clk ) begin
        s798_val_n7 <= s797_val_n7;
    end
    always @(posedge \clk ) begin
        \s799_val  <= \s798_val ;
    end
    always @(posedge \clk ) begin
        s799_val_n1 <= s798_val_n1;
    end
    always @(posedge \clk ) begin
        s799_val_n2 <= s798_val_n2;
    end
    always @(posedge \clk ) begin
        s799_val_n3 <= s798_val_n3;
    end
    always @(posedge \clk ) begin
        s799_val_n4 <= s798_val_n4;
    end
    always @(posedge \clk ) begin
        s799_val_n5 <= s798_val_n5;
    end
    always @(posedge \clk ) begin
        s799_val_n6 <= s798_val_n6;
    end
    always @(posedge \clk ) begin
        s799_val_n7 <= s798_val_n7;
    end
    always @(posedge \clk ) begin
        \s800_val  <= \s799_val ;
    end
    always @(posedge \clk ) begin
        s800_val_n1 <= s799_val_n1;
    end
    always @(posedge \clk ) begin
        s800_val_n2 <= s799_val_n2;
    end
    always @(posedge \clk ) begin
        s800_val_n3 <= s799_val_n3;
    end
    always @(posedge \clk ) begin
        s800_val_n4 <= s799_val_n4;
    end
    always @(posedge \clk ) begin
        s800_val_n5 <= s799_val_n5;
    end
    always @(posedge \clk ) begin
        s800_val_n6 <= s799_val_n6;
    end
    always @(posedge \clk ) begin
        s800_val_n7 <= s799_val_n7;
    end
    always @(posedge \clk ) begin
        \s801_val  <= \s800_val ;
    end
    always @(posedge \clk ) begin
        s801_val_n1 <= s800_val_n1;
    end
    always @(posedge \clk ) begin
        s801_val_n2 <= s800_val_n2;
    end
    always @(posedge \clk ) begin
        s801_val_n3 <= s800_val_n3;
    end
    always @(posedge \clk ) begin
        s801_val_n4 <= s800_val_n4;
    end
    always @(posedge \clk ) begin
        s801_val_n5 <= s800_val_n5;
    end
    always @(posedge \clk ) begin
        s801_val_n6 <= s800_val_n6;
    end
    always @(posedge \clk ) begin
        s801_val_n7 <= s800_val_n7;
    end
    always @(posedge \clk ) begin
        s801_val_n8 <= val_n8;
    end
    always @(posedge \clk ) begin
        \s802_val  <= \s801_val ;
    end
    always @(posedge \clk ) begin
        s802_val_n1 <= s801_val_n1;
    end
    always @(posedge \clk ) begin
        s802_val_n2 <= s801_val_n2;
    end
    always @(posedge \clk ) begin
        s802_val_n3 <= s801_val_n3;
    end
    always @(posedge \clk ) begin
        s802_val_n4 <= s801_val_n4;
    end
    always @(posedge \clk ) begin
        s802_val_n5 <= s801_val_n5;
    end
    always @(posedge \clk ) begin
        s802_val_n6 <= s801_val_n6;
    end
    always @(posedge \clk ) begin
        s802_val_n7 <= s801_val_n7;
    end
    always @(posedge \clk ) begin
        s802_val_n8 <= s801_val_n8;
    end
    always @(posedge \clk ) begin
        \s803_val  <= \s802_val ;
    end
    always @(posedge \clk ) begin
        s803_val_n1 <= s802_val_n1;
    end
    always @(posedge \clk ) begin
        s803_val_n2 <= s802_val_n2;
    end
    always @(posedge \clk ) begin
        s803_val_n3 <= s802_val_n3;
    end
    always @(posedge \clk ) begin
        s803_val_n4 <= s802_val_n4;
    end
    always @(posedge \clk ) begin
        s803_val_n5 <= s802_val_n5;
    end
    always @(posedge \clk ) begin
        s803_val_n6 <= s802_val_n6;
    end
    always @(posedge \clk ) begin
        s803_val_n7 <= s802_val_n7;
    end
    always @(posedge \clk ) begin
        s803_val_n8 <= s802_val_n8;
    end
    always @(posedge \clk ) begin
        \s804_val  <= \s803_val ;
    end
    always @(posedge \clk ) begin
        s804_val_n1 <= s803_val_n1;
    end
    always @(posedge \clk ) begin
        s804_val_n2 <= s803_val_n2;
    end
    always @(posedge \clk ) begin
        s804_val_n3 <= s803_val_n3;
    end
    always @(posedge \clk ) begin
        s804_val_n4 <= s803_val_n4;
    end
    always @(posedge \clk ) begin
        s804_val_n5 <= s803_val_n5;
    end
    always @(posedge \clk ) begin
        s804_val_n6 <= s803_val_n6;
    end
    always @(posedge \clk ) begin
        s804_val_n7 <= s803_val_n7;
    end
    always @(posedge \clk ) begin
        s804_val_n8 <= s803_val_n8;
    end
    always @(posedge \clk ) begin
        \s805_val  <= \s804_val ;
    end
    always @(posedge \clk ) begin
        s805_val_n1 <= s804_val_n1;
    end
    always @(posedge \clk ) begin
        s805_val_n2 <= s804_val_n2;
    end
    always @(posedge \clk ) begin
        s805_val_n3 <= s804_val_n3;
    end
    always @(posedge \clk ) begin
        s805_val_n4 <= s804_val_n4;
    end
    always @(posedge \clk ) begin
        s805_val_n5 <= s804_val_n5;
    end
    always @(posedge \clk ) begin
        s805_val_n6 <= s804_val_n6;
    end
    always @(posedge \clk ) begin
        s805_val_n7 <= s804_val_n7;
    end
    always @(posedge \clk ) begin
        s805_val_n8 <= s804_val_n8;
    end
    always @(posedge \clk ) begin
        \s806_val  <= \s805_val ;
    end
    always @(posedge \clk ) begin
        s806_val_n1 <= s805_val_n1;
    end
    always @(posedge \clk ) begin
        s806_val_n2 <= s805_val_n2;
    end
    always @(posedge \clk ) begin
        s806_val_n3 <= s805_val_n3;
    end
    always @(posedge \clk ) begin
        s806_val_n4 <= s805_val_n4;
    end
    always @(posedge \clk ) begin
        s806_val_n5 <= s805_val_n5;
    end
    always @(posedge \clk ) begin
        s806_val_n6 <= s805_val_n6;
    end
    always @(posedge \clk ) begin
        s806_val_n7 <= s805_val_n7;
    end
    always @(posedge \clk ) begin
        s806_val_n8 <= s805_val_n8;
    end
    always @(posedge \clk ) begin
        \s807_val  <= \s806_val ;
    end
    always @(posedge \clk ) begin
        s807_val_n1 <= s806_val_n1;
    end
    always @(posedge \clk ) begin
        s807_val_n2 <= s806_val_n2;
    end
    always @(posedge \clk ) begin
        s807_val_n3 <= s806_val_n3;
    end
    always @(posedge \clk ) begin
        s807_val_n4 <= s806_val_n4;
    end
    always @(posedge \clk ) begin
        s807_val_n5 <= s806_val_n5;
    end
    always @(posedge \clk ) begin
        s807_val_n6 <= s806_val_n6;
    end
    always @(posedge \clk ) begin
        s807_val_n7 <= s806_val_n7;
    end
    always @(posedge \clk ) begin
        s807_val_n8 <= s806_val_n8;
    end
    always @(posedge \clk ) begin
        \s808_val  <= \s807_val ;
    end
    always @(posedge \clk ) begin
        s808_val_n1 <= s807_val_n1;
    end
    always @(posedge \clk ) begin
        s808_val_n2 <= s807_val_n2;
    end
    always @(posedge \clk ) begin
        s808_val_n3 <= s807_val_n3;
    end
    always @(posedge \clk ) begin
        s808_val_n4 <= s807_val_n4;
    end
    always @(posedge \clk ) begin
        s808_val_n5 <= s807_val_n5;
    end
    always @(posedge \clk ) begin
        s808_val_n6 <= s807_val_n6;
    end
    always @(posedge \clk ) begin
        s808_val_n7 <= s807_val_n7;
    end
    always @(posedge \clk ) begin
        s808_val_n8 <= s807_val_n8;
    end
    always @(posedge \clk ) begin
        \s809_val  <= \s808_val ;
    end
    always @(posedge \clk ) begin
        s809_val_n1 <= s808_val_n1;
    end
    always @(posedge \clk ) begin
        s809_val_n2 <= s808_val_n2;
    end
    always @(posedge \clk ) begin
        s809_val_n3 <= s808_val_n3;
    end
    always @(posedge \clk ) begin
        s809_val_n4 <= s808_val_n4;
    end
    always @(posedge \clk ) begin
        s809_val_n5 <= s808_val_n5;
    end
    always @(posedge \clk ) begin
        s809_val_n6 <= s808_val_n6;
    end
    always @(posedge \clk ) begin
        s809_val_n7 <= s808_val_n7;
    end
    always @(posedge \clk ) begin
        s809_val_n8 <= s808_val_n8;
    end
    always @(posedge \clk ) begin
        \s810_val  <= \s809_val ;
    end
    always @(posedge \clk ) begin
        s810_val_n1 <= s809_val_n1;
    end
    always @(posedge \clk ) begin
        s810_val_n2 <= s809_val_n2;
    end
    always @(posedge \clk ) begin
        s810_val_n3 <= s809_val_n3;
    end
    always @(posedge \clk ) begin
        s810_val_n4 <= s809_val_n4;
    end
    always @(posedge \clk ) begin
        s810_val_n5 <= s809_val_n5;
    end
    always @(posedge \clk ) begin
        s810_val_n6 <= s809_val_n6;
    end
    always @(posedge \clk ) begin
        s810_val_n7 <= s809_val_n7;
    end
    always @(posedge \clk ) begin
        s810_val_n8 <= s809_val_n8;
    end
    always @(posedge \clk ) begin
        \s811_val  <= \s810_val ;
    end
    always @(posedge \clk ) begin
        s811_val_n1 <= s810_val_n1;
    end
    always @(posedge \clk ) begin
        s811_val_n2 <= s810_val_n2;
    end
    always @(posedge \clk ) begin
        s811_val_n3 <= s810_val_n3;
    end
    always @(posedge \clk ) begin
        s811_val_n4 <= s810_val_n4;
    end
    always @(posedge \clk ) begin
        s811_val_n5 <= s810_val_n5;
    end
    always @(posedge \clk ) begin
        s811_val_n6 <= s810_val_n6;
    end
    always @(posedge \clk ) begin
        s811_val_n7 <= s810_val_n7;
    end
    always @(posedge \clk ) begin
        s811_val_n8 <= s810_val_n8;
    end
    always @(posedge \clk ) begin
        \s812_val  <= \s811_val ;
    end
    always @(posedge \clk ) begin
        s812_val_n1 <= s811_val_n1;
    end
    always @(posedge \clk ) begin
        s812_val_n2 <= s811_val_n2;
    end
    always @(posedge \clk ) begin
        s812_val_n3 <= s811_val_n3;
    end
    always @(posedge \clk ) begin
        s812_val_n4 <= s811_val_n4;
    end
    always @(posedge \clk ) begin
        s812_val_n5 <= s811_val_n5;
    end
    always @(posedge \clk ) begin
        s812_val_n6 <= s811_val_n6;
    end
    always @(posedge \clk ) begin
        s812_val_n7 <= s811_val_n7;
    end
    always @(posedge \clk ) begin
        s812_val_n8 <= s811_val_n8;
    end
    always @(posedge \clk ) begin
        \s813_val  <= \s812_val ;
    end
    always @(posedge \clk ) begin
        s813_val_n1 <= s812_val_n1;
    end
    always @(posedge \clk ) begin
        s813_val_n2 <= s812_val_n2;
    end
    always @(posedge \clk ) begin
        s813_val_n3 <= s812_val_n3;
    end
    always @(posedge \clk ) begin
        s813_val_n4 <= s812_val_n4;
    end
    always @(posedge \clk ) begin
        s813_val_n5 <= s812_val_n5;
    end
    always @(posedge \clk ) begin
        s813_val_n6 <= s812_val_n6;
    end
    always @(posedge \clk ) begin
        s813_val_n7 <= s812_val_n7;
    end
    always @(posedge \clk ) begin
        s813_val_n8 <= s812_val_n8;
    end
    always @(posedge \clk ) begin
        \s814_val  <= \s813_val ;
    end
    always @(posedge \clk ) begin
        s814_val_n1 <= s813_val_n1;
    end
    always @(posedge \clk ) begin
        s814_val_n2 <= s813_val_n2;
    end
    always @(posedge \clk ) begin
        s814_val_n3 <= s813_val_n3;
    end
    always @(posedge \clk ) begin
        s814_val_n4 <= s813_val_n4;
    end
    always @(posedge \clk ) begin
        s814_val_n5 <= s813_val_n5;
    end
    always @(posedge \clk ) begin
        s814_val_n6 <= s813_val_n6;
    end
    always @(posedge \clk ) begin
        s814_val_n7 <= s813_val_n7;
    end
    always @(posedge \clk ) begin
        s814_val_n8 <= s813_val_n8;
    end
    always @(posedge \clk ) begin
        \s815_val  <= \s814_val ;
    end
    always @(posedge \clk ) begin
        s815_val_n1 <= s814_val_n1;
    end
    always @(posedge \clk ) begin
        s815_val_n2 <= s814_val_n2;
    end
    always @(posedge \clk ) begin
        s815_val_n3 <= s814_val_n3;
    end
    always @(posedge \clk ) begin
        s815_val_n4 <= s814_val_n4;
    end
    always @(posedge \clk ) begin
        s815_val_n5 <= s814_val_n5;
    end
    always @(posedge \clk ) begin
        s815_val_n6 <= s814_val_n6;
    end
    always @(posedge \clk ) begin
        s815_val_n7 <= s814_val_n7;
    end
    always @(posedge \clk ) begin
        s815_val_n8 <= s814_val_n8;
    end
    always @(posedge \clk ) begin
        \s816_val  <= \s815_val ;
    end
    always @(posedge \clk ) begin
        s816_val_n1 <= s815_val_n1;
    end
    always @(posedge \clk ) begin
        s816_val_n2 <= s815_val_n2;
    end
    always @(posedge \clk ) begin
        s816_val_n3 <= s815_val_n3;
    end
    always @(posedge \clk ) begin
        s816_val_n4 <= s815_val_n4;
    end
    always @(posedge \clk ) begin
        s816_val_n5 <= s815_val_n5;
    end
    always @(posedge \clk ) begin
        s816_val_n6 <= s815_val_n6;
    end
    always @(posedge \clk ) begin
        s816_val_n7 <= s815_val_n7;
    end
    always @(posedge \clk ) begin
        s816_val_n8 <= s815_val_n8;
    end
    always @(posedge \clk ) begin
        \s817_val  <= \s816_val ;
    end
    always @(posedge \clk ) begin
        s817_val_n1 <= s816_val_n1;
    end
    always @(posedge \clk ) begin
        s817_val_n2 <= s816_val_n2;
    end
    always @(posedge \clk ) begin
        s817_val_n3 <= s816_val_n3;
    end
    always @(posedge \clk ) begin
        s817_val_n4 <= s816_val_n4;
    end
    always @(posedge \clk ) begin
        s817_val_n5 <= s816_val_n5;
    end
    always @(posedge \clk ) begin
        s817_val_n6 <= s816_val_n6;
    end
    always @(posedge \clk ) begin
        s817_val_n7 <= s816_val_n7;
    end
    always @(posedge \clk ) begin
        s817_val_n8 <= s816_val_n8;
    end
    always @(posedge \clk ) begin
        \s818_val  <= \s817_val ;
    end
    always @(posedge \clk ) begin
        s818_val_n1 <= s817_val_n1;
    end
    always @(posedge \clk ) begin
        s818_val_n2 <= s817_val_n2;
    end
    always @(posedge \clk ) begin
        s818_val_n3 <= s817_val_n3;
    end
    always @(posedge \clk ) begin
        s818_val_n4 <= s817_val_n4;
    end
    always @(posedge \clk ) begin
        s818_val_n5 <= s817_val_n5;
    end
    always @(posedge \clk ) begin
        s818_val_n6 <= s817_val_n6;
    end
    always @(posedge \clk ) begin
        s818_val_n7 <= s817_val_n7;
    end
    always @(posedge \clk ) begin
        s818_val_n8 <= s817_val_n8;
    end
    always @(posedge \clk ) begin
        \s819_val  <= \s818_val ;
    end
    always @(posedge \clk ) begin
        s819_val_n1 <= s818_val_n1;
    end
    always @(posedge \clk ) begin
        s819_val_n2 <= s818_val_n2;
    end
    always @(posedge \clk ) begin
        s819_val_n3 <= s818_val_n3;
    end
    always @(posedge \clk ) begin
        s819_val_n4 <= s818_val_n4;
    end
    always @(posedge \clk ) begin
        s819_val_n5 <= s818_val_n5;
    end
    always @(posedge \clk ) begin
        s819_val_n6 <= s818_val_n6;
    end
    always @(posedge \clk ) begin
        s819_val_n7 <= s818_val_n7;
    end
    always @(posedge \clk ) begin
        s819_val_n8 <= s818_val_n8;
    end
    always @(posedge \clk ) begin
        \s820_val  <= \s819_val ;
    end
    always @(posedge \clk ) begin
        s820_val_n1 <= s819_val_n1;
    end
    always @(posedge \clk ) begin
        s820_val_n2 <= s819_val_n2;
    end
    always @(posedge \clk ) begin
        s820_val_n3 <= s819_val_n3;
    end
    always @(posedge \clk ) begin
        s820_val_n4 <= s819_val_n4;
    end
    always @(posedge \clk ) begin
        s820_val_n5 <= s819_val_n5;
    end
    always @(posedge \clk ) begin
        s820_val_n6 <= s819_val_n6;
    end
    always @(posedge \clk ) begin
        s820_val_n7 <= s819_val_n7;
    end
    always @(posedge \clk ) begin
        s820_val_n8 <= s819_val_n8;
    end
    always @(posedge \clk ) begin
        \s821_val  <= \s820_val ;
    end
    always @(posedge \clk ) begin
        s821_val_n1 <= s820_val_n1;
    end
    always @(posedge \clk ) begin
        s821_val_n2 <= s820_val_n2;
    end
    always @(posedge \clk ) begin
        s821_val_n3 <= s820_val_n3;
    end
    always @(posedge \clk ) begin
        s821_val_n4 <= s820_val_n4;
    end
    always @(posedge \clk ) begin
        s821_val_n5 <= s820_val_n5;
    end
    always @(posedge \clk ) begin
        s821_val_n6 <= s820_val_n6;
    end
    always @(posedge \clk ) begin
        s821_val_n7 <= s820_val_n7;
    end
    always @(posedge \clk ) begin
        s821_val_n8 <= s820_val_n8;
    end
    always @(posedge \clk ) begin
        \s822_val  <= \s821_val ;
    end
    always @(posedge \clk ) begin
        s822_val_n1 <= s821_val_n1;
    end
    always @(posedge \clk ) begin
        s822_val_n2 <= s821_val_n2;
    end
    always @(posedge \clk ) begin
        s822_val_n3 <= s821_val_n3;
    end
    always @(posedge \clk ) begin
        s822_val_n4 <= s821_val_n4;
    end
    always @(posedge \clk ) begin
        s822_val_n5 <= s821_val_n5;
    end
    always @(posedge \clk ) begin
        s822_val_n6 <= s821_val_n6;
    end
    always @(posedge \clk ) begin
        s822_val_n7 <= s821_val_n7;
    end
    always @(posedge \clk ) begin
        s822_val_n8 <= s821_val_n8;
    end
    always @(posedge \clk ) begin
        \s823_val  <= \s822_val ;
    end
    always @(posedge \clk ) begin
        s823_val_n1 <= s822_val_n1;
    end
    always @(posedge \clk ) begin
        s823_val_n2 <= s822_val_n2;
    end
    always @(posedge \clk ) begin
        s823_val_n3 <= s822_val_n3;
    end
    always @(posedge \clk ) begin
        s823_val_n4 <= s822_val_n4;
    end
    always @(posedge \clk ) begin
        s823_val_n5 <= s822_val_n5;
    end
    always @(posedge \clk ) begin
        s823_val_n6 <= s822_val_n6;
    end
    always @(posedge \clk ) begin
        s823_val_n7 <= s822_val_n7;
    end
    always @(posedge \clk ) begin
        s823_val_n8 <= s822_val_n8;
    end
    always @(posedge \clk ) begin
        \s824_val  <= \s823_val ;
    end
    always @(posedge \clk ) begin
        s824_val_n1 <= s823_val_n1;
    end
    always @(posedge \clk ) begin
        s824_val_n2 <= s823_val_n2;
    end
    always @(posedge \clk ) begin
        s824_val_n3 <= s823_val_n3;
    end
    always @(posedge \clk ) begin
        s824_val_n4 <= s823_val_n4;
    end
    always @(posedge \clk ) begin
        s824_val_n5 <= s823_val_n5;
    end
    always @(posedge \clk ) begin
        s824_val_n6 <= s823_val_n6;
    end
    always @(posedge \clk ) begin
        s824_val_n7 <= s823_val_n7;
    end
    always @(posedge \clk ) begin
        s824_val_n8 <= s823_val_n8;
    end
    always @(posedge \clk ) begin
        \s825_val  <= \s824_val ;
    end
    always @(posedge \clk ) begin
        s825_val_n1 <= s824_val_n1;
    end
    always @(posedge \clk ) begin
        s825_val_n2 <= s824_val_n2;
    end
    always @(posedge \clk ) begin
        s825_val_n3 <= s824_val_n3;
    end
    always @(posedge \clk ) begin
        s825_val_n4 <= s824_val_n4;
    end
    always @(posedge \clk ) begin
        s825_val_n5 <= s824_val_n5;
    end
    always @(posedge \clk ) begin
        s825_val_n6 <= s824_val_n6;
    end
    always @(posedge \clk ) begin
        s825_val_n7 <= s824_val_n7;
    end
    always @(posedge \clk ) begin
        s825_val_n8 <= s824_val_n8;
    end
    always @(posedge \clk ) begin
        \s826_val  <= \s825_val ;
    end
    always @(posedge \clk ) begin
        s826_val_n1 <= s825_val_n1;
    end
    always @(posedge \clk ) begin
        s826_val_n2 <= s825_val_n2;
    end
    always @(posedge \clk ) begin
        s826_val_n3 <= s825_val_n3;
    end
    always @(posedge \clk ) begin
        s826_val_n4 <= s825_val_n4;
    end
    always @(posedge \clk ) begin
        s826_val_n5 <= s825_val_n5;
    end
    always @(posedge \clk ) begin
        s826_val_n6 <= s825_val_n6;
    end
    always @(posedge \clk ) begin
        s826_val_n7 <= s825_val_n7;
    end
    always @(posedge \clk ) begin
        s826_val_n8 <= s825_val_n8;
    end
    always @(posedge \clk ) begin
        \s827_val  <= \s826_val ;
    end
    always @(posedge \clk ) begin
        s827_val_n1 <= s826_val_n1;
    end
    always @(posedge \clk ) begin
        s827_val_n2 <= s826_val_n2;
    end
    always @(posedge \clk ) begin
        s827_val_n3 <= s826_val_n3;
    end
    always @(posedge \clk ) begin
        s827_val_n4 <= s826_val_n4;
    end
    always @(posedge \clk ) begin
        s827_val_n5 <= s826_val_n5;
    end
    always @(posedge \clk ) begin
        s827_val_n6 <= s826_val_n6;
    end
    always @(posedge \clk ) begin
        s827_val_n7 <= s826_val_n7;
    end
    always @(posedge \clk ) begin
        s827_val_n8 <= s826_val_n8;
    end
    always @(posedge \clk ) begin
        \s828_val  <= \s827_val ;
    end
    always @(posedge \clk ) begin
        s828_val_n1 <= s827_val_n1;
    end
    always @(posedge \clk ) begin
        s828_val_n2 <= s827_val_n2;
    end
    always @(posedge \clk ) begin
        s828_val_n3 <= s827_val_n3;
    end
    always @(posedge \clk ) begin
        s828_val_n4 <= s827_val_n4;
    end
    always @(posedge \clk ) begin
        s828_val_n5 <= s827_val_n5;
    end
    always @(posedge \clk ) begin
        s828_val_n6 <= s827_val_n6;
    end
    always @(posedge \clk ) begin
        s828_val_n7 <= s827_val_n7;
    end
    always @(posedge \clk ) begin
        s828_val_n8 <= s827_val_n8;
    end
    always @(posedge \clk ) begin
        \s829_val  <= \s828_val ;
    end
    always @(posedge \clk ) begin
        s829_val_n1 <= s828_val_n1;
    end
    always @(posedge \clk ) begin
        s829_val_n2 <= s828_val_n2;
    end
    always @(posedge \clk ) begin
        s829_val_n3 <= s828_val_n3;
    end
    always @(posedge \clk ) begin
        s829_val_n4 <= s828_val_n4;
    end
    always @(posedge \clk ) begin
        s829_val_n5 <= s828_val_n5;
    end
    always @(posedge \clk ) begin
        s829_val_n6 <= s828_val_n6;
    end
    always @(posedge \clk ) begin
        s829_val_n7 <= s828_val_n7;
    end
    always @(posedge \clk ) begin
        s829_val_n8 <= s828_val_n8;
    end
    always @(posedge \clk ) begin
        \s830_val  <= \s829_val ;
    end
    always @(posedge \clk ) begin
        s830_val_n1 <= s829_val_n1;
    end
    always @(posedge \clk ) begin
        s830_val_n2 <= s829_val_n2;
    end
    always @(posedge \clk ) begin
        s830_val_n3 <= s829_val_n3;
    end
    always @(posedge \clk ) begin
        s830_val_n4 <= s829_val_n4;
    end
    always @(posedge \clk ) begin
        s830_val_n5 <= s829_val_n5;
    end
    always @(posedge \clk ) begin
        s830_val_n6 <= s829_val_n6;
    end
    always @(posedge \clk ) begin
        s830_val_n7 <= s829_val_n7;
    end
    always @(posedge \clk ) begin
        s830_val_n8 <= s829_val_n8;
    end
    always @(posedge \clk ) begin
        \s831_val  <= \s830_val ;
    end
    always @(posedge \clk ) begin
        s831_val_n1 <= s830_val_n1;
    end
    always @(posedge \clk ) begin
        s831_val_n2 <= s830_val_n2;
    end
    always @(posedge \clk ) begin
        s831_val_n3 <= s830_val_n3;
    end
    always @(posedge \clk ) begin
        s831_val_n4 <= s830_val_n4;
    end
    always @(posedge \clk ) begin
        s831_val_n5 <= s830_val_n5;
    end
    always @(posedge \clk ) begin
        s831_val_n6 <= s830_val_n6;
    end
    always @(posedge \clk ) begin
        s831_val_n7 <= s830_val_n7;
    end
    always @(posedge \clk ) begin
        s831_val_n8 <= s830_val_n8;
    end
    always @(posedge \clk ) begin
        \s832_val  <= \s831_val ;
    end
    always @(posedge \clk ) begin
        s832_val_n1 <= s831_val_n1;
    end
    always @(posedge \clk ) begin
        s832_val_n2 <= s831_val_n2;
    end
    always @(posedge \clk ) begin
        s832_val_n3 <= s831_val_n3;
    end
    always @(posedge \clk ) begin
        s832_val_n4 <= s831_val_n4;
    end
    always @(posedge \clk ) begin
        s832_val_n5 <= s831_val_n5;
    end
    always @(posedge \clk ) begin
        s832_val_n6 <= s831_val_n6;
    end
    always @(posedge \clk ) begin
        s832_val_n7 <= s831_val_n7;
    end
    always @(posedge \clk ) begin
        s832_val_n8 <= s831_val_n8;
    end
    always @(posedge \clk ) begin
        \s833_val  <= \s832_val ;
    end
    always @(posedge \clk ) begin
        s833_val_n1 <= s832_val_n1;
    end
    always @(posedge \clk ) begin
        s833_val_n2 <= s832_val_n2;
    end
    always @(posedge \clk ) begin
        s833_val_n3 <= s832_val_n3;
    end
    always @(posedge \clk ) begin
        s833_val_n4 <= s832_val_n4;
    end
    always @(posedge \clk ) begin
        s833_val_n5 <= s832_val_n5;
    end
    always @(posedge \clk ) begin
        s833_val_n6 <= s832_val_n6;
    end
    always @(posedge \clk ) begin
        s833_val_n7 <= s832_val_n7;
    end
    always @(posedge \clk ) begin
        s833_val_n8 <= s832_val_n8;
    end
    always @(posedge \clk ) begin
        \s834_val  <= \s833_val ;
    end
    always @(posedge \clk ) begin
        s834_val_n1 <= s833_val_n1;
    end
    always @(posedge \clk ) begin
        s834_val_n2 <= s833_val_n2;
    end
    always @(posedge \clk ) begin
        s834_val_n3 <= s833_val_n3;
    end
    always @(posedge \clk ) begin
        s834_val_n4 <= s833_val_n4;
    end
    always @(posedge \clk ) begin
        s834_val_n5 <= s833_val_n5;
    end
    always @(posedge \clk ) begin
        s834_val_n6 <= s833_val_n6;
    end
    always @(posedge \clk ) begin
        s834_val_n7 <= s833_val_n7;
    end
    always @(posedge \clk ) begin
        s834_val_n8 <= s833_val_n8;
    end
    always @(posedge \clk ) begin
        \s835_val  <= \s834_val ;
    end
    always @(posedge \clk ) begin
        s835_val_n1 <= s834_val_n1;
    end
    always @(posedge \clk ) begin
        s835_val_n2 <= s834_val_n2;
    end
    always @(posedge \clk ) begin
        s835_val_n3 <= s834_val_n3;
    end
    always @(posedge \clk ) begin
        s835_val_n4 <= s834_val_n4;
    end
    always @(posedge \clk ) begin
        s835_val_n5 <= s834_val_n5;
    end
    always @(posedge \clk ) begin
        s835_val_n6 <= s834_val_n6;
    end
    always @(posedge \clk ) begin
        s835_val_n7 <= s834_val_n7;
    end
    always @(posedge \clk ) begin
        s835_val_n8 <= s834_val_n8;
    end
    always @(posedge \clk ) begin
        \s836_val  <= \s835_val ;
    end
    always @(posedge \clk ) begin
        s836_val_n1 <= s835_val_n1;
    end
    always @(posedge \clk ) begin
        s836_val_n2 <= s835_val_n2;
    end
    always @(posedge \clk ) begin
        s836_val_n3 <= s835_val_n3;
    end
    always @(posedge \clk ) begin
        s836_val_n4 <= s835_val_n4;
    end
    always @(posedge \clk ) begin
        s836_val_n5 <= s835_val_n5;
    end
    always @(posedge \clk ) begin
        s836_val_n6 <= s835_val_n6;
    end
    always @(posedge \clk ) begin
        s836_val_n7 <= s835_val_n7;
    end
    always @(posedge \clk ) begin
        s836_val_n8 <= s835_val_n8;
    end
    always @(posedge \clk ) begin
        \s837_val  <= \s836_val ;
    end
    always @(posedge \clk ) begin
        s837_val_n1 <= s836_val_n1;
    end
    always @(posedge \clk ) begin
        s837_val_n2 <= s836_val_n2;
    end
    always @(posedge \clk ) begin
        s837_val_n3 <= s836_val_n3;
    end
    always @(posedge \clk ) begin
        s837_val_n4 <= s836_val_n4;
    end
    always @(posedge \clk ) begin
        s837_val_n5 <= s836_val_n5;
    end
    always @(posedge \clk ) begin
        s837_val_n6 <= s836_val_n6;
    end
    always @(posedge \clk ) begin
        s837_val_n7 <= s836_val_n7;
    end
    always @(posedge \clk ) begin
        s837_val_n8 <= s836_val_n8;
    end
    always @(posedge \clk ) begin
        \s838_val  <= \s837_val ;
    end
    always @(posedge \clk ) begin
        s838_val_n1 <= s837_val_n1;
    end
    always @(posedge \clk ) begin
        s838_val_n2 <= s837_val_n2;
    end
    always @(posedge \clk ) begin
        s838_val_n3 <= s837_val_n3;
    end
    always @(posedge \clk ) begin
        s838_val_n4 <= s837_val_n4;
    end
    always @(posedge \clk ) begin
        s838_val_n5 <= s837_val_n5;
    end
    always @(posedge \clk ) begin
        s838_val_n6 <= s837_val_n6;
    end
    always @(posedge \clk ) begin
        s838_val_n7 <= s837_val_n7;
    end
    always @(posedge \clk ) begin
        s838_val_n8 <= s837_val_n8;
    end
    always @(posedge \clk ) begin
        \s839_val  <= \s838_val ;
    end
    always @(posedge \clk ) begin
        s839_val_n1 <= s838_val_n1;
    end
    always @(posedge \clk ) begin
        s839_val_n2 <= s838_val_n2;
    end
    always @(posedge \clk ) begin
        s839_val_n3 <= s838_val_n3;
    end
    always @(posedge \clk ) begin
        s839_val_n4 <= s838_val_n4;
    end
    always @(posedge \clk ) begin
        s839_val_n5 <= s838_val_n5;
    end
    always @(posedge \clk ) begin
        s839_val_n6 <= s838_val_n6;
    end
    always @(posedge \clk ) begin
        s839_val_n7 <= s838_val_n7;
    end
    always @(posedge \clk ) begin
        s839_val_n8 <= s838_val_n8;
    end
    always @(posedge \clk ) begin
        \s840_val  <= \s839_val ;
    end
    always @(posedge \clk ) begin
        s840_val_n1 <= s839_val_n1;
    end
    always @(posedge \clk ) begin
        s840_val_n2 <= s839_val_n2;
    end
    always @(posedge \clk ) begin
        s840_val_n3 <= s839_val_n3;
    end
    always @(posedge \clk ) begin
        s840_val_n4 <= s839_val_n4;
    end
    always @(posedge \clk ) begin
        s840_val_n5 <= s839_val_n5;
    end
    always @(posedge \clk ) begin
        s840_val_n6 <= s839_val_n6;
    end
    always @(posedge \clk ) begin
        s840_val_n7 <= s839_val_n7;
    end
    always @(posedge \clk ) begin
        s840_val_n8 <= s839_val_n8;
    end
    always @(posedge \clk ) begin
        \s841_val  <= \s840_val ;
    end
    always @(posedge \clk ) begin
        s841_val_n1 <= s840_val_n1;
    end
    always @(posedge \clk ) begin
        s841_val_n2 <= s840_val_n2;
    end
    always @(posedge \clk ) begin
        s841_val_n3 <= s840_val_n3;
    end
    always @(posedge \clk ) begin
        s841_val_n4 <= s840_val_n4;
    end
    always @(posedge \clk ) begin
        s841_val_n5 <= s840_val_n5;
    end
    always @(posedge \clk ) begin
        s841_val_n6 <= s840_val_n6;
    end
    always @(posedge \clk ) begin
        s841_val_n7 <= s840_val_n7;
    end
    always @(posedge \clk ) begin
        s841_val_n8 <= s840_val_n8;
    end
    always @(posedge \clk ) begin
        \s842_val  <= \s841_val ;
    end
    always @(posedge \clk ) begin
        s842_val_n1 <= s841_val_n1;
    end
    always @(posedge \clk ) begin
        s842_val_n2 <= s841_val_n2;
    end
    always @(posedge \clk ) begin
        s842_val_n3 <= s841_val_n3;
    end
    always @(posedge \clk ) begin
        s842_val_n4 <= s841_val_n4;
    end
    always @(posedge \clk ) begin
        s842_val_n5 <= s841_val_n5;
    end
    always @(posedge \clk ) begin
        s842_val_n6 <= s841_val_n6;
    end
    always @(posedge \clk ) begin
        s842_val_n7 <= s841_val_n7;
    end
    always @(posedge \clk ) begin
        s842_val_n8 <= s841_val_n8;
    end
    always @(posedge \clk ) begin
        \s843_val  <= \s842_val ;
    end
    always @(posedge \clk ) begin
        s843_val_n1 <= s842_val_n1;
    end
    always @(posedge \clk ) begin
        s843_val_n2 <= s842_val_n2;
    end
    always @(posedge \clk ) begin
        s843_val_n3 <= s842_val_n3;
    end
    always @(posedge \clk ) begin
        s843_val_n4 <= s842_val_n4;
    end
    always @(posedge \clk ) begin
        s843_val_n5 <= s842_val_n5;
    end
    always @(posedge \clk ) begin
        s843_val_n6 <= s842_val_n6;
    end
    always @(posedge \clk ) begin
        s843_val_n7 <= s842_val_n7;
    end
    always @(posedge \clk ) begin
        s843_val_n8 <= s842_val_n8;
    end
    always @(posedge \clk ) begin
        \s844_val  <= \s843_val ;
    end
    always @(posedge \clk ) begin
        s844_val_n1 <= s843_val_n1;
    end
    always @(posedge \clk ) begin
        s844_val_n2 <= s843_val_n2;
    end
    always @(posedge \clk ) begin
        s844_val_n3 <= s843_val_n3;
    end
    always @(posedge \clk ) begin
        s844_val_n4 <= s843_val_n4;
    end
    always @(posedge \clk ) begin
        s844_val_n5 <= s843_val_n5;
    end
    always @(posedge \clk ) begin
        s844_val_n6 <= s843_val_n6;
    end
    always @(posedge \clk ) begin
        s844_val_n7 <= s843_val_n7;
    end
    always @(posedge \clk ) begin
        s844_val_n8 <= s843_val_n8;
    end
    always @(posedge \clk ) begin
        \s845_val  <= \s844_val ;
    end
    always @(posedge \clk ) begin
        s845_val_n1 <= s844_val_n1;
    end
    always @(posedge \clk ) begin
        s845_val_n2 <= s844_val_n2;
    end
    always @(posedge \clk ) begin
        s845_val_n3 <= s844_val_n3;
    end
    always @(posedge \clk ) begin
        s845_val_n4 <= s844_val_n4;
    end
    always @(posedge \clk ) begin
        s845_val_n5 <= s844_val_n5;
    end
    always @(posedge \clk ) begin
        s845_val_n6 <= s844_val_n6;
    end
    always @(posedge \clk ) begin
        s845_val_n7 <= s844_val_n7;
    end
    always @(posedge \clk ) begin
        s845_val_n8 <= s844_val_n8;
    end
    always @(posedge \clk ) begin
        \s846_val  <= \s845_val ;
    end
    always @(posedge \clk ) begin
        s846_val_n1 <= s845_val_n1;
    end
    always @(posedge \clk ) begin
        s846_val_n2 <= s845_val_n2;
    end
    always @(posedge \clk ) begin
        s846_val_n3 <= s845_val_n3;
    end
    always @(posedge \clk ) begin
        s846_val_n4 <= s845_val_n4;
    end
    always @(posedge \clk ) begin
        s846_val_n5 <= s845_val_n5;
    end
    always @(posedge \clk ) begin
        s846_val_n6 <= s845_val_n6;
    end
    always @(posedge \clk ) begin
        s846_val_n7 <= s845_val_n7;
    end
    always @(posedge \clk ) begin
        s846_val_n8 <= s845_val_n8;
    end
    always @(posedge \clk ) begin
        \s847_val  <= \s846_val ;
    end
    always @(posedge \clk ) begin
        s847_val_n1 <= s846_val_n1;
    end
    always @(posedge \clk ) begin
        s847_val_n2 <= s846_val_n2;
    end
    always @(posedge \clk ) begin
        s847_val_n3 <= s846_val_n3;
    end
    always @(posedge \clk ) begin
        s847_val_n4 <= s846_val_n4;
    end
    always @(posedge \clk ) begin
        s847_val_n5 <= s846_val_n5;
    end
    always @(posedge \clk ) begin
        s847_val_n6 <= s846_val_n6;
    end
    always @(posedge \clk ) begin
        s847_val_n7 <= s846_val_n7;
    end
    always @(posedge \clk ) begin
        s847_val_n8 <= s846_val_n8;
    end
    always @(posedge \clk ) begin
        \s848_val  <= \s847_val ;
    end
    always @(posedge \clk ) begin
        s848_val_n1 <= s847_val_n1;
    end
    always @(posedge \clk ) begin
        s848_val_n2 <= s847_val_n2;
    end
    always @(posedge \clk ) begin
        s848_val_n3 <= s847_val_n3;
    end
    always @(posedge \clk ) begin
        s848_val_n4 <= s847_val_n4;
    end
    always @(posedge \clk ) begin
        s848_val_n5 <= s847_val_n5;
    end
    always @(posedge \clk ) begin
        s848_val_n6 <= s847_val_n6;
    end
    always @(posedge \clk ) begin
        s848_val_n7 <= s847_val_n7;
    end
    always @(posedge \clk ) begin
        s848_val_n8 <= s847_val_n8;
    end
    always @(posedge \clk ) begin
        \s849_val  <= \s848_val ;
    end
    always @(posedge \clk ) begin
        s849_val_n1 <= s848_val_n1;
    end
    always @(posedge \clk ) begin
        s849_val_n2 <= s848_val_n2;
    end
    always @(posedge \clk ) begin
        s849_val_n3 <= s848_val_n3;
    end
    always @(posedge \clk ) begin
        s849_val_n4 <= s848_val_n4;
    end
    always @(posedge \clk ) begin
        s849_val_n5 <= s848_val_n5;
    end
    always @(posedge \clk ) begin
        s849_val_n6 <= s848_val_n6;
    end
    always @(posedge \clk ) begin
        s849_val_n7 <= s848_val_n7;
    end
    always @(posedge \clk ) begin
        s849_val_n8 <= s848_val_n8;
    end
    always @(posedge \clk ) begin
        \s850_val  <= \s849_val ;
    end
    always @(posedge \clk ) begin
        s850_val_n1 <= s849_val_n1;
    end
    always @(posedge \clk ) begin
        s850_val_n2 <= s849_val_n2;
    end
    always @(posedge \clk ) begin
        s850_val_n3 <= s849_val_n3;
    end
    always @(posedge \clk ) begin
        s850_val_n4 <= s849_val_n4;
    end
    always @(posedge \clk ) begin
        s850_val_n5 <= s849_val_n5;
    end
    always @(posedge \clk ) begin
        s850_val_n6 <= s849_val_n6;
    end
    always @(posedge \clk ) begin
        s850_val_n7 <= s849_val_n7;
    end
    always @(posedge \clk ) begin
        s850_val_n8 <= s849_val_n8;
    end
    always @(posedge \clk ) begin
        \s851_val  <= \s850_val ;
    end
    always @(posedge \clk ) begin
        s851_val_n1 <= s850_val_n1;
    end
    always @(posedge \clk ) begin
        s851_val_n2 <= s850_val_n2;
    end
    always @(posedge \clk ) begin
        s851_val_n3 <= s850_val_n3;
    end
    always @(posedge \clk ) begin
        s851_val_n4 <= s850_val_n4;
    end
    always @(posedge \clk ) begin
        s851_val_n5 <= s850_val_n5;
    end
    always @(posedge \clk ) begin
        s851_val_n6 <= s850_val_n6;
    end
    always @(posedge \clk ) begin
        s851_val_n7 <= s850_val_n7;
    end
    always @(posedge \clk ) begin
        s851_val_n8 <= s850_val_n8;
    end
    always @(posedge \clk ) begin
        \s852_val  <= \s851_val ;
    end
    always @(posedge \clk ) begin
        s852_val_n1 <= s851_val_n1;
    end
    always @(posedge \clk ) begin
        s852_val_n2 <= s851_val_n2;
    end
    always @(posedge \clk ) begin
        s852_val_n3 <= s851_val_n3;
    end
    always @(posedge \clk ) begin
        s852_val_n4 <= s851_val_n4;
    end
    always @(posedge \clk ) begin
        s852_val_n5 <= s851_val_n5;
    end
    always @(posedge \clk ) begin
        s852_val_n6 <= s851_val_n6;
    end
    always @(posedge \clk ) begin
        s852_val_n7 <= s851_val_n7;
    end
    always @(posedge \clk ) begin
        s852_val_n8 <= s851_val_n8;
    end
    always @(posedge \clk ) begin
        \s853_val  <= \s852_val ;
    end
    always @(posedge \clk ) begin
        s853_val_n1 <= s852_val_n1;
    end
    always @(posedge \clk ) begin
        s853_val_n2 <= s852_val_n2;
    end
    always @(posedge \clk ) begin
        s853_val_n3 <= s852_val_n3;
    end
    always @(posedge \clk ) begin
        s853_val_n4 <= s852_val_n4;
    end
    always @(posedge \clk ) begin
        s853_val_n5 <= s852_val_n5;
    end
    always @(posedge \clk ) begin
        s853_val_n6 <= s852_val_n6;
    end
    always @(posedge \clk ) begin
        s853_val_n7 <= s852_val_n7;
    end
    always @(posedge \clk ) begin
        s853_val_n8 <= s852_val_n8;
    end
    always @(posedge \clk ) begin
        \s854_val  <= \s853_val ;
    end
    always @(posedge \clk ) begin
        s854_val_n1 <= s853_val_n1;
    end
    always @(posedge \clk ) begin
        s854_val_n2 <= s853_val_n2;
    end
    always @(posedge \clk ) begin
        s854_val_n3 <= s853_val_n3;
    end
    always @(posedge \clk ) begin
        s854_val_n4 <= s853_val_n4;
    end
    always @(posedge \clk ) begin
        s854_val_n5 <= s853_val_n5;
    end
    always @(posedge \clk ) begin
        s854_val_n6 <= s853_val_n6;
    end
    always @(posedge \clk ) begin
        s854_val_n7 <= s853_val_n7;
    end
    always @(posedge \clk ) begin
        s854_val_n8 <= s853_val_n8;
    end
    always @(posedge \clk ) begin
        \s855_val  <= \s854_val ;
    end
    always @(posedge \clk ) begin
        s855_val_n1 <= s854_val_n1;
    end
    always @(posedge \clk ) begin
        s855_val_n2 <= s854_val_n2;
    end
    always @(posedge \clk ) begin
        s855_val_n3 <= s854_val_n3;
    end
    always @(posedge \clk ) begin
        s855_val_n4 <= s854_val_n4;
    end
    always @(posedge \clk ) begin
        s855_val_n5 <= s854_val_n5;
    end
    always @(posedge \clk ) begin
        s855_val_n6 <= s854_val_n6;
    end
    always @(posedge \clk ) begin
        s855_val_n7 <= s854_val_n7;
    end
    always @(posedge \clk ) begin
        s855_val_n8 <= s854_val_n8;
    end
    always @(posedge \clk ) begin
        \s856_val  <= \s855_val ;
    end
    always @(posedge \clk ) begin
        s856_val_n1 <= s855_val_n1;
    end
    always @(posedge \clk ) begin
        s856_val_n2 <= s855_val_n2;
    end
    always @(posedge \clk ) begin
        s856_val_n3 <= s855_val_n3;
    end
    always @(posedge \clk ) begin
        s856_val_n4 <= s855_val_n4;
    end
    always @(posedge \clk ) begin
        s856_val_n5 <= s855_val_n5;
    end
    always @(posedge \clk ) begin
        s856_val_n6 <= s855_val_n6;
    end
    always @(posedge \clk ) begin
        s856_val_n7 <= s855_val_n7;
    end
    always @(posedge \clk ) begin
        s856_val_n8 <= s855_val_n8;
    end
    always @(posedge \clk ) begin
        \s857_val  <= \s856_val ;
    end
    always @(posedge \clk ) begin
        s857_val_n1 <= s856_val_n1;
    end
    always @(posedge \clk ) begin
        s857_val_n2 <= s856_val_n2;
    end
    always @(posedge \clk ) begin
        s857_val_n3 <= s856_val_n3;
    end
    always @(posedge \clk ) begin
        s857_val_n4 <= s856_val_n4;
    end
    always @(posedge \clk ) begin
        s857_val_n5 <= s856_val_n5;
    end
    always @(posedge \clk ) begin
        s857_val_n6 <= s856_val_n6;
    end
    always @(posedge \clk ) begin
        s857_val_n7 <= s856_val_n7;
    end
    always @(posedge \clk ) begin
        s857_val_n8 <= s856_val_n8;
    end
    always @(posedge \clk ) begin
        \s858_val  <= \s857_val ;
    end
    always @(posedge \clk ) begin
        s858_val_n1 <= s857_val_n1;
    end
    always @(posedge \clk ) begin
        s858_val_n2 <= s857_val_n2;
    end
    always @(posedge \clk ) begin
        s858_val_n3 <= s857_val_n3;
    end
    always @(posedge \clk ) begin
        s858_val_n4 <= s857_val_n4;
    end
    always @(posedge \clk ) begin
        s858_val_n5 <= s857_val_n5;
    end
    always @(posedge \clk ) begin
        s858_val_n6 <= s857_val_n6;
    end
    always @(posedge \clk ) begin
        s858_val_n7 <= s857_val_n7;
    end
    always @(posedge \clk ) begin
        s858_val_n8 <= s857_val_n8;
    end
    always @(posedge \clk ) begin
        \s859_val  <= \s858_val ;
    end
    always @(posedge \clk ) begin
        s859_val_n1 <= s858_val_n1;
    end
    always @(posedge \clk ) begin
        s859_val_n2 <= s858_val_n2;
    end
    always @(posedge \clk ) begin
        s859_val_n3 <= s858_val_n3;
    end
    always @(posedge \clk ) begin
        s859_val_n4 <= s858_val_n4;
    end
    always @(posedge \clk ) begin
        s859_val_n5 <= s858_val_n5;
    end
    always @(posedge \clk ) begin
        s859_val_n6 <= s858_val_n6;
    end
    always @(posedge \clk ) begin
        s859_val_n7 <= s858_val_n7;
    end
    always @(posedge \clk ) begin
        s859_val_n8 <= s858_val_n8;
    end
    always @(posedge \clk ) begin
        \s860_val  <= \s859_val ;
    end
    always @(posedge \clk ) begin
        s860_val_n1 <= s859_val_n1;
    end
    always @(posedge \clk ) begin
        s860_val_n2 <= s859_val_n2;
    end
    always @(posedge \clk ) begin
        s860_val_n3 <= s859_val_n3;
    end
    always @(posedge \clk ) begin
        s860_val_n4 <= s859_val_n4;
    end
    always @(posedge \clk ) begin
        s860_val_n5 <= s859_val_n5;
    end
    always @(posedge \clk ) begin
        s860_val_n6 <= s859_val_n6;
    end
    always @(posedge \clk ) begin
        s860_val_n7 <= s859_val_n7;
    end
    always @(posedge \clk ) begin
        s860_val_n8 <= s859_val_n8;
    end
    always @(posedge \clk ) begin
        \s861_val  <= \s860_val ;
    end
    always @(posedge \clk ) begin
        s861_val_n1 <= s860_val_n1;
    end
    always @(posedge \clk ) begin
        s861_val_n2 <= s860_val_n2;
    end
    always @(posedge \clk ) begin
        s861_val_n3 <= s860_val_n3;
    end
    always @(posedge \clk ) begin
        s861_val_n4 <= s860_val_n4;
    end
    always @(posedge \clk ) begin
        s861_val_n5 <= s860_val_n5;
    end
    always @(posedge \clk ) begin
        s861_val_n6 <= s860_val_n6;
    end
    always @(posedge \clk ) begin
        s861_val_n7 <= s860_val_n7;
    end
    always @(posedge \clk ) begin
        s861_val_n8 <= s860_val_n8;
    end
    always @(posedge \clk ) begin
        \s862_val  <= \s861_val ;
    end
    always @(posedge \clk ) begin
        s862_val_n1 <= s861_val_n1;
    end
    always @(posedge \clk ) begin
        s862_val_n2 <= s861_val_n2;
    end
    always @(posedge \clk ) begin
        s862_val_n3 <= s861_val_n3;
    end
    always @(posedge \clk ) begin
        s862_val_n4 <= s861_val_n4;
    end
    always @(posedge \clk ) begin
        s862_val_n5 <= s861_val_n5;
    end
    always @(posedge \clk ) begin
        s862_val_n6 <= s861_val_n6;
    end
    always @(posedge \clk ) begin
        s862_val_n7 <= s861_val_n7;
    end
    always @(posedge \clk ) begin
        s862_val_n8 <= s861_val_n8;
    end
    always @(posedge \clk ) begin
        \s863_val  <= \s862_val ;
    end
    always @(posedge \clk ) begin
        s863_val_n1 <= s862_val_n1;
    end
    always @(posedge \clk ) begin
        s863_val_n2 <= s862_val_n2;
    end
    always @(posedge \clk ) begin
        s863_val_n3 <= s862_val_n3;
    end
    always @(posedge \clk ) begin
        s863_val_n4 <= s862_val_n4;
    end
    always @(posedge \clk ) begin
        s863_val_n5 <= s862_val_n5;
    end
    always @(posedge \clk ) begin
        s863_val_n6 <= s862_val_n6;
    end
    always @(posedge \clk ) begin
        s863_val_n7 <= s862_val_n7;
    end
    always @(posedge \clk ) begin
        s863_val_n8 <= s862_val_n8;
    end
    always @(posedge \clk ) begin
        \s864_val  <= \s863_val ;
    end
    always @(posedge \clk ) begin
        s864_val_n1 <= s863_val_n1;
    end
    always @(posedge \clk ) begin
        s864_val_n2 <= s863_val_n2;
    end
    always @(posedge \clk ) begin
        s864_val_n3 <= s863_val_n3;
    end
    always @(posedge \clk ) begin
        s864_val_n4 <= s863_val_n4;
    end
    always @(posedge \clk ) begin
        s864_val_n5 <= s863_val_n5;
    end
    always @(posedge \clk ) begin
        s864_val_n6 <= s863_val_n6;
    end
    always @(posedge \clk ) begin
        s864_val_n7 <= s863_val_n7;
    end
    always @(posedge \clk ) begin
        s864_val_n8 <= s863_val_n8;
    end
    always @(posedge \clk ) begin
        \s865_val  <= \s864_val ;
    end
    always @(posedge \clk ) begin
        s865_val_n1 <= s864_val_n1;
    end
    always @(posedge \clk ) begin
        s865_val_n2 <= s864_val_n2;
    end
    always @(posedge \clk ) begin
        s865_val_n3 <= s864_val_n3;
    end
    always @(posedge \clk ) begin
        s865_val_n4 <= s864_val_n4;
    end
    always @(posedge \clk ) begin
        s865_val_n5 <= s864_val_n5;
    end
    always @(posedge \clk ) begin
        s865_val_n6 <= s864_val_n6;
    end
    always @(posedge \clk ) begin
        s865_val_n7 <= s864_val_n7;
    end
    always @(posedge \clk ) begin
        s865_val_n8 <= s864_val_n8;
    end
    always @(posedge \clk ) begin
        \s866_val  <= \s865_val ;
    end
    always @(posedge \clk ) begin
        s866_val_n1 <= s865_val_n1;
    end
    always @(posedge \clk ) begin
        s866_val_n2 <= s865_val_n2;
    end
    always @(posedge \clk ) begin
        s866_val_n3 <= s865_val_n3;
    end
    always @(posedge \clk ) begin
        s866_val_n4 <= s865_val_n4;
    end
    always @(posedge \clk ) begin
        s866_val_n5 <= s865_val_n5;
    end
    always @(posedge \clk ) begin
        s866_val_n6 <= s865_val_n6;
    end
    always @(posedge \clk ) begin
        s866_val_n7 <= s865_val_n7;
    end
    always @(posedge \clk ) begin
        s866_val_n8 <= s865_val_n8;
    end
    always @(posedge \clk ) begin
        \s867_val  <= \s866_val ;
    end
    always @(posedge \clk ) begin
        s867_val_n1 <= s866_val_n1;
    end
    always @(posedge \clk ) begin
        s867_val_n2 <= s866_val_n2;
    end
    always @(posedge \clk ) begin
        s867_val_n3 <= s866_val_n3;
    end
    always @(posedge \clk ) begin
        s867_val_n4 <= s866_val_n4;
    end
    always @(posedge \clk ) begin
        s867_val_n5 <= s866_val_n5;
    end
    always @(posedge \clk ) begin
        s867_val_n6 <= s866_val_n6;
    end
    always @(posedge \clk ) begin
        s867_val_n7 <= s866_val_n7;
    end
    always @(posedge \clk ) begin
        s867_val_n8 <= s866_val_n8;
    end
    always @(posedge \clk ) begin
        \s868_val  <= \s867_val ;
    end
    always @(posedge \clk ) begin
        s868_val_n1 <= s867_val_n1;
    end
    always @(posedge \clk ) begin
        s868_val_n2 <= s867_val_n2;
    end
    always @(posedge \clk ) begin
        s868_val_n3 <= s867_val_n3;
    end
    always @(posedge \clk ) begin
        s868_val_n4 <= s867_val_n4;
    end
    always @(posedge \clk ) begin
        s868_val_n5 <= s867_val_n5;
    end
    always @(posedge \clk ) begin
        s868_val_n6 <= s867_val_n6;
    end
    always @(posedge \clk ) begin
        s868_val_n7 <= s867_val_n7;
    end
    always @(posedge \clk ) begin
        s868_val_n8 <= s867_val_n8;
    end
    always @(posedge \clk ) begin
        \s869_val  <= \s868_val ;
    end
    always @(posedge \clk ) begin
        s869_val_n1 <= s868_val_n1;
    end
    always @(posedge \clk ) begin
        s869_val_n2 <= s868_val_n2;
    end
    always @(posedge \clk ) begin
        s869_val_n3 <= s868_val_n3;
    end
    always @(posedge \clk ) begin
        s869_val_n4 <= s868_val_n4;
    end
    always @(posedge \clk ) begin
        s869_val_n5 <= s868_val_n5;
    end
    always @(posedge \clk ) begin
        s869_val_n6 <= s868_val_n6;
    end
    always @(posedge \clk ) begin
        s869_val_n7 <= s868_val_n7;
    end
    always @(posedge \clk ) begin
        s869_val_n8 <= s868_val_n8;
    end
    always @(posedge \clk ) begin
        \s870_val  <= \s869_val ;
    end
    always @(posedge \clk ) begin
        s870_val_n1 <= s869_val_n1;
    end
    always @(posedge \clk ) begin
        s870_val_n2 <= s869_val_n2;
    end
    always @(posedge \clk ) begin
        s870_val_n3 <= s869_val_n3;
    end
    always @(posedge \clk ) begin
        s870_val_n4 <= s869_val_n4;
    end
    always @(posedge \clk ) begin
        s870_val_n5 <= s869_val_n5;
    end
    always @(posedge \clk ) begin
        s870_val_n6 <= s869_val_n6;
    end
    always @(posedge \clk ) begin
        s870_val_n7 <= s869_val_n7;
    end
    always @(posedge \clk ) begin
        s870_val_n8 <= s869_val_n8;
    end
    always @(posedge \clk ) begin
        \s871_val  <= \s870_val ;
    end
    always @(posedge \clk ) begin
        s871_val_n1 <= s870_val_n1;
    end
    always @(posedge \clk ) begin
        s871_val_n2 <= s870_val_n2;
    end
    always @(posedge \clk ) begin
        s871_val_n3 <= s870_val_n3;
    end
    always @(posedge \clk ) begin
        s871_val_n4 <= s870_val_n4;
    end
    always @(posedge \clk ) begin
        s871_val_n5 <= s870_val_n5;
    end
    always @(posedge \clk ) begin
        s871_val_n6 <= s870_val_n6;
    end
    always @(posedge \clk ) begin
        s871_val_n7 <= s870_val_n7;
    end
    always @(posedge \clk ) begin
        s871_val_n8 <= s870_val_n8;
    end
    always @(posedge \clk ) begin
        \s872_val  <= \s871_val ;
    end
    always @(posedge \clk ) begin
        s872_val_n1 <= s871_val_n1;
    end
    always @(posedge \clk ) begin
        s872_val_n2 <= s871_val_n2;
    end
    always @(posedge \clk ) begin
        s872_val_n3 <= s871_val_n3;
    end
    always @(posedge \clk ) begin
        s872_val_n4 <= s871_val_n4;
    end
    always @(posedge \clk ) begin
        s872_val_n5 <= s871_val_n5;
    end
    always @(posedge \clk ) begin
        s872_val_n6 <= s871_val_n6;
    end
    always @(posedge \clk ) begin
        s872_val_n7 <= s871_val_n7;
    end
    always @(posedge \clk ) begin
        s872_val_n8 <= s871_val_n8;
    end
    always @(posedge \clk ) begin
        \s873_val  <= \s872_val ;
    end
    always @(posedge \clk ) begin
        s873_val_n1 <= s872_val_n1;
    end
    always @(posedge \clk ) begin
        s873_val_n2 <= s872_val_n2;
    end
    always @(posedge \clk ) begin
        s873_val_n3 <= s872_val_n3;
    end
    always @(posedge \clk ) begin
        s873_val_n4 <= s872_val_n4;
    end
    always @(posedge \clk ) begin
        s873_val_n5 <= s872_val_n5;
    end
    always @(posedge \clk ) begin
        s873_val_n6 <= s872_val_n6;
    end
    always @(posedge \clk ) begin
        s873_val_n7 <= s872_val_n7;
    end
    always @(posedge \clk ) begin
        s873_val_n8 <= s872_val_n8;
    end
    always @(posedge \clk ) begin
        \s874_val  <= \s873_val ;
    end
    always @(posedge \clk ) begin
        s874_val_n1 <= s873_val_n1;
    end
    always @(posedge \clk ) begin
        s874_val_n2 <= s873_val_n2;
    end
    always @(posedge \clk ) begin
        s874_val_n3 <= s873_val_n3;
    end
    always @(posedge \clk ) begin
        s874_val_n4 <= s873_val_n4;
    end
    always @(posedge \clk ) begin
        s874_val_n5 <= s873_val_n5;
    end
    always @(posedge \clk ) begin
        s874_val_n6 <= s873_val_n6;
    end
    always @(posedge \clk ) begin
        s874_val_n7 <= s873_val_n7;
    end
    always @(posedge \clk ) begin
        s874_val_n8 <= s873_val_n8;
    end
    always @(posedge \clk ) begin
        \s875_val  <= \s874_val ;
    end
    always @(posedge \clk ) begin
        s875_val_n1 <= s874_val_n1;
    end
    always @(posedge \clk ) begin
        s875_val_n2 <= s874_val_n2;
    end
    always @(posedge \clk ) begin
        s875_val_n3 <= s874_val_n3;
    end
    always @(posedge \clk ) begin
        s875_val_n4 <= s874_val_n4;
    end
    always @(posedge \clk ) begin
        s875_val_n5 <= s874_val_n5;
    end
    always @(posedge \clk ) begin
        s875_val_n6 <= s874_val_n6;
    end
    always @(posedge \clk ) begin
        s875_val_n7 <= s874_val_n7;
    end
    always @(posedge \clk ) begin
        s875_val_n8 <= s874_val_n8;
    end
    always @(posedge \clk ) begin
        \s876_val  <= \s875_val ;
    end
    always @(posedge \clk ) begin
        s876_val_n1 <= s875_val_n1;
    end
    always @(posedge \clk ) begin
        s876_val_n2 <= s875_val_n2;
    end
    always @(posedge \clk ) begin
        s876_val_n3 <= s875_val_n3;
    end
    always @(posedge \clk ) begin
        s876_val_n4 <= s875_val_n4;
    end
    always @(posedge \clk ) begin
        s876_val_n5 <= s875_val_n5;
    end
    always @(posedge \clk ) begin
        s876_val_n6 <= s875_val_n6;
    end
    always @(posedge \clk ) begin
        s876_val_n7 <= s875_val_n7;
    end
    always @(posedge \clk ) begin
        s876_val_n8 <= s875_val_n8;
    end
    always @(posedge \clk ) begin
        \s877_val  <= \s876_val ;
    end
    always @(posedge \clk ) begin
        s877_val_n1 <= s876_val_n1;
    end
    always @(posedge \clk ) begin
        s877_val_n2 <= s876_val_n2;
    end
    always @(posedge \clk ) begin
        s877_val_n3 <= s876_val_n3;
    end
    always @(posedge \clk ) begin
        s877_val_n4 <= s876_val_n4;
    end
    always @(posedge \clk ) begin
        s877_val_n5 <= s876_val_n5;
    end
    always @(posedge \clk ) begin
        s877_val_n6 <= s876_val_n6;
    end
    always @(posedge \clk ) begin
        s877_val_n7 <= s876_val_n7;
    end
    always @(posedge \clk ) begin
        s877_val_n8 <= s876_val_n8;
    end
    always @(posedge \clk ) begin
        \s878_val  <= \s877_val ;
    end
    always @(posedge \clk ) begin
        s878_val_n1 <= s877_val_n1;
    end
    always @(posedge \clk ) begin
        s878_val_n2 <= s877_val_n2;
    end
    always @(posedge \clk ) begin
        s878_val_n3 <= s877_val_n3;
    end
    always @(posedge \clk ) begin
        s878_val_n4 <= s877_val_n4;
    end
    always @(posedge \clk ) begin
        s878_val_n5 <= s877_val_n5;
    end
    always @(posedge \clk ) begin
        s878_val_n6 <= s877_val_n6;
    end
    always @(posedge \clk ) begin
        s878_val_n7 <= s877_val_n7;
    end
    always @(posedge \clk ) begin
        s878_val_n8 <= s877_val_n8;
    end
    always @(posedge \clk ) begin
        \s879_val  <= \s878_val ;
    end
    always @(posedge \clk ) begin
        s879_val_n1 <= s878_val_n1;
    end
    always @(posedge \clk ) begin
        s879_val_n2 <= s878_val_n2;
    end
    always @(posedge \clk ) begin
        s879_val_n3 <= s878_val_n3;
    end
    always @(posedge \clk ) begin
        s879_val_n4 <= s878_val_n4;
    end
    always @(posedge \clk ) begin
        s879_val_n5 <= s878_val_n5;
    end
    always @(posedge \clk ) begin
        s879_val_n6 <= s878_val_n6;
    end
    always @(posedge \clk ) begin
        s879_val_n7 <= s878_val_n7;
    end
    always @(posedge \clk ) begin
        s879_val_n8 <= s878_val_n8;
    end
    always @(posedge \clk ) begin
        \s880_val  <= \s879_val ;
    end
    always @(posedge \clk ) begin
        s880_val_n1 <= s879_val_n1;
    end
    always @(posedge \clk ) begin
        s880_val_n2 <= s879_val_n2;
    end
    always @(posedge \clk ) begin
        s880_val_n3 <= s879_val_n3;
    end
    always @(posedge \clk ) begin
        s880_val_n4 <= s879_val_n4;
    end
    always @(posedge \clk ) begin
        s880_val_n5 <= s879_val_n5;
    end
    always @(posedge \clk ) begin
        s880_val_n6 <= s879_val_n6;
    end
    always @(posedge \clk ) begin
        s880_val_n7 <= s879_val_n7;
    end
    always @(posedge \clk ) begin
        s880_val_n8 <= s879_val_n8;
    end
    always @(posedge \clk ) begin
        \s881_val  <= \s880_val ;
    end
    always @(posedge \clk ) begin
        s881_val_n1 <= s880_val_n1;
    end
    always @(posedge \clk ) begin
        s881_val_n2 <= s880_val_n2;
    end
    always @(posedge \clk ) begin
        s881_val_n3 <= s880_val_n3;
    end
    always @(posedge \clk ) begin
        s881_val_n4 <= s880_val_n4;
    end
    always @(posedge \clk ) begin
        s881_val_n5 <= s880_val_n5;
    end
    always @(posedge \clk ) begin
        s881_val_n6 <= s880_val_n6;
    end
    always @(posedge \clk ) begin
        s881_val_n7 <= s880_val_n7;
    end
    always @(posedge \clk ) begin
        s881_val_n8 <= s880_val_n8;
    end
    always @(posedge \clk ) begin
        \s882_val  <= \s881_val ;
    end
    always @(posedge \clk ) begin
        s882_val_n1 <= s881_val_n1;
    end
    always @(posedge \clk ) begin
        s882_val_n2 <= s881_val_n2;
    end
    always @(posedge \clk ) begin
        s882_val_n3 <= s881_val_n3;
    end
    always @(posedge \clk ) begin
        s882_val_n4 <= s881_val_n4;
    end
    always @(posedge \clk ) begin
        s882_val_n5 <= s881_val_n5;
    end
    always @(posedge \clk ) begin
        s882_val_n6 <= s881_val_n6;
    end
    always @(posedge \clk ) begin
        s882_val_n7 <= s881_val_n7;
    end
    always @(posedge \clk ) begin
        s882_val_n8 <= s881_val_n8;
    end
    always @(posedge \clk ) begin
        \s883_val  <= \s882_val ;
    end
    always @(posedge \clk ) begin
        s883_val_n1 <= s882_val_n1;
    end
    always @(posedge \clk ) begin
        s883_val_n2 <= s882_val_n2;
    end
    always @(posedge \clk ) begin
        s883_val_n3 <= s882_val_n3;
    end
    always @(posedge \clk ) begin
        s883_val_n4 <= s882_val_n4;
    end
    always @(posedge \clk ) begin
        s883_val_n5 <= s882_val_n5;
    end
    always @(posedge \clk ) begin
        s883_val_n6 <= s882_val_n6;
    end
    always @(posedge \clk ) begin
        s883_val_n7 <= s882_val_n7;
    end
    always @(posedge \clk ) begin
        s883_val_n8 <= s882_val_n8;
    end
    always @(posedge \clk ) begin
        \s884_val  <= \s883_val ;
    end
    always @(posedge \clk ) begin
        s884_val_n1 <= s883_val_n1;
    end
    always @(posedge \clk ) begin
        s884_val_n2 <= s883_val_n2;
    end
    always @(posedge \clk ) begin
        s884_val_n3 <= s883_val_n3;
    end
    always @(posedge \clk ) begin
        s884_val_n4 <= s883_val_n4;
    end
    always @(posedge \clk ) begin
        s884_val_n5 <= s883_val_n5;
    end
    always @(posedge \clk ) begin
        s884_val_n6 <= s883_val_n6;
    end
    always @(posedge \clk ) begin
        s884_val_n7 <= s883_val_n7;
    end
    always @(posedge \clk ) begin
        s884_val_n8 <= s883_val_n8;
    end
    always @(posedge \clk ) begin
        \s885_val  <= \s884_val ;
    end
    always @(posedge \clk ) begin
        s885_val_n1 <= s884_val_n1;
    end
    always @(posedge \clk ) begin
        s885_val_n2 <= s884_val_n2;
    end
    always @(posedge \clk ) begin
        s885_val_n3 <= s884_val_n3;
    end
    always @(posedge \clk ) begin
        s885_val_n4 <= s884_val_n4;
    end
    always @(posedge \clk ) begin
        s885_val_n5 <= s884_val_n5;
    end
    always @(posedge \clk ) begin
        s885_val_n6 <= s884_val_n6;
    end
    always @(posedge \clk ) begin
        s885_val_n7 <= s884_val_n7;
    end
    always @(posedge \clk ) begin
        s885_val_n8 <= s884_val_n8;
    end
    always @(posedge \clk ) begin
        \s886_val  <= \s885_val ;
    end
    always @(posedge \clk ) begin
        s886_val_n1 <= s885_val_n1;
    end
    always @(posedge \clk ) begin
        s886_val_n2 <= s885_val_n2;
    end
    always @(posedge \clk ) begin
        s886_val_n3 <= s885_val_n3;
    end
    always @(posedge \clk ) begin
        s886_val_n4 <= s885_val_n4;
    end
    always @(posedge \clk ) begin
        s886_val_n5 <= s885_val_n5;
    end
    always @(posedge \clk ) begin
        s886_val_n6 <= s885_val_n6;
    end
    always @(posedge \clk ) begin
        s886_val_n7 <= s885_val_n7;
    end
    always @(posedge \clk ) begin
        s886_val_n8 <= s885_val_n8;
    end
    always @(posedge \clk ) begin
        \s887_val  <= \s886_val ;
    end
    always @(posedge \clk ) begin
        s887_val_n1 <= s886_val_n1;
    end
    always @(posedge \clk ) begin
        s887_val_n2 <= s886_val_n2;
    end
    always @(posedge \clk ) begin
        s887_val_n3 <= s886_val_n3;
    end
    always @(posedge \clk ) begin
        s887_val_n4 <= s886_val_n4;
    end
    always @(posedge \clk ) begin
        s887_val_n5 <= s886_val_n5;
    end
    always @(posedge \clk ) begin
        s887_val_n6 <= s886_val_n6;
    end
    always @(posedge \clk ) begin
        s887_val_n7 <= s886_val_n7;
    end
    always @(posedge \clk ) begin
        s887_val_n8 <= s886_val_n8;
    end
    always @(posedge \clk ) begin
        \s888_val  <= \s887_val ;
    end
    always @(posedge \clk ) begin
        s888_val_n1 <= s887_val_n1;
    end
    always @(posedge \clk ) begin
        s888_val_n2 <= s887_val_n2;
    end
    always @(posedge \clk ) begin
        s888_val_n3 <= s887_val_n3;
    end
    always @(posedge \clk ) begin
        s888_val_n4 <= s887_val_n4;
    end
    always @(posedge \clk ) begin
        s888_val_n5 <= s887_val_n5;
    end
    always @(posedge \clk ) begin
        s888_val_n6 <= s887_val_n6;
    end
    always @(posedge \clk ) begin
        s888_val_n7 <= s887_val_n7;
    end
    always @(posedge \clk ) begin
        s888_val_n8 <= s887_val_n8;
    end
    always @(posedge \clk ) begin
        \s889_val  <= \s888_val ;
    end
    always @(posedge \clk ) begin
        s889_val_n1 <= s888_val_n1;
    end
    always @(posedge \clk ) begin
        s889_val_n2 <= s888_val_n2;
    end
    always @(posedge \clk ) begin
        s889_val_n3 <= s888_val_n3;
    end
    always @(posedge \clk ) begin
        s889_val_n4 <= s888_val_n4;
    end
    always @(posedge \clk ) begin
        s889_val_n5 <= s888_val_n5;
    end
    always @(posedge \clk ) begin
        s889_val_n6 <= s888_val_n6;
    end
    always @(posedge \clk ) begin
        s889_val_n7 <= s888_val_n7;
    end
    always @(posedge \clk ) begin
        s889_val_n8 <= s888_val_n8;
    end
    always @(posedge \clk ) begin
        \s890_val  <= \s889_val ;
    end
    always @(posedge \clk ) begin
        s890_val_n1 <= s889_val_n1;
    end
    always @(posedge \clk ) begin
        s890_val_n2 <= s889_val_n2;
    end
    always @(posedge \clk ) begin
        s890_val_n3 <= s889_val_n3;
    end
    always @(posedge \clk ) begin
        s890_val_n4 <= s889_val_n4;
    end
    always @(posedge \clk ) begin
        s890_val_n5 <= s889_val_n5;
    end
    always @(posedge \clk ) begin
        s890_val_n6 <= s889_val_n6;
    end
    always @(posedge \clk ) begin
        s890_val_n7 <= s889_val_n7;
    end
    always @(posedge \clk ) begin
        s890_val_n8 <= s889_val_n8;
    end
    always @(posedge \clk ) begin
        \s891_val  <= \s890_val ;
    end
    always @(posedge \clk ) begin
        s891_val_n1 <= s890_val_n1;
    end
    always @(posedge \clk ) begin
        s891_val_n2 <= s890_val_n2;
    end
    always @(posedge \clk ) begin
        s891_val_n3 <= s890_val_n3;
    end
    always @(posedge \clk ) begin
        s891_val_n4 <= s890_val_n4;
    end
    always @(posedge \clk ) begin
        s891_val_n5 <= s890_val_n5;
    end
    always @(posedge \clk ) begin
        s891_val_n6 <= s890_val_n6;
    end
    always @(posedge \clk ) begin
        s891_val_n7 <= s890_val_n7;
    end
    always @(posedge \clk ) begin
        s891_val_n8 <= s890_val_n8;
    end
    always @(posedge \clk ) begin
        \s892_val  <= \s891_val ;
    end
    always @(posedge \clk ) begin
        s892_val_n1 <= s891_val_n1;
    end
    always @(posedge \clk ) begin
        s892_val_n2 <= s891_val_n2;
    end
    always @(posedge \clk ) begin
        s892_val_n3 <= s891_val_n3;
    end
    always @(posedge \clk ) begin
        s892_val_n4 <= s891_val_n4;
    end
    always @(posedge \clk ) begin
        s892_val_n5 <= s891_val_n5;
    end
    always @(posedge \clk ) begin
        s892_val_n6 <= s891_val_n6;
    end
    always @(posedge \clk ) begin
        s892_val_n7 <= s891_val_n7;
    end
    always @(posedge \clk ) begin
        s892_val_n8 <= s891_val_n8;
    end
    always @(posedge \clk ) begin
        \s893_val  <= \s892_val ;
    end
    always @(posedge \clk ) begin
        s893_val_n1 <= s892_val_n1;
    end
    always @(posedge \clk ) begin
        s893_val_n2 <= s892_val_n2;
    end
    always @(posedge \clk ) begin
        s893_val_n3 <= s892_val_n3;
    end
    always @(posedge \clk ) begin
        s893_val_n4 <= s892_val_n4;
    end
    always @(posedge \clk ) begin
        s893_val_n5 <= s892_val_n5;
    end
    always @(posedge \clk ) begin
        s893_val_n6 <= s892_val_n6;
    end
    always @(posedge \clk ) begin
        s893_val_n7 <= s892_val_n7;
    end
    always @(posedge \clk ) begin
        s893_val_n8 <= s892_val_n8;
    end
    always @(posedge \clk ) begin
        \s894_val  <= \s893_val ;
    end
    always @(posedge \clk ) begin
        s894_val_n1 <= s893_val_n1;
    end
    always @(posedge \clk ) begin
        s894_val_n2 <= s893_val_n2;
    end
    always @(posedge \clk ) begin
        s894_val_n3 <= s893_val_n3;
    end
    always @(posedge \clk ) begin
        s894_val_n4 <= s893_val_n4;
    end
    always @(posedge \clk ) begin
        s894_val_n5 <= s893_val_n5;
    end
    always @(posedge \clk ) begin
        s894_val_n6 <= s893_val_n6;
    end
    always @(posedge \clk ) begin
        s894_val_n7 <= s893_val_n7;
    end
    always @(posedge \clk ) begin
        s894_val_n8 <= s893_val_n8;
    end
    always @(posedge \clk ) begin
        \s895_val  <= \s894_val ;
    end
    always @(posedge \clk ) begin
        s895_val_n1 <= s894_val_n1;
    end
    always @(posedge \clk ) begin
        s895_val_n2 <= s894_val_n2;
    end
    always @(posedge \clk ) begin
        s895_val_n3 <= s894_val_n3;
    end
    always @(posedge \clk ) begin
        s895_val_n4 <= s894_val_n4;
    end
    always @(posedge \clk ) begin
        s895_val_n5 <= s894_val_n5;
    end
    always @(posedge \clk ) begin
        s895_val_n6 <= s894_val_n6;
    end
    always @(posedge \clk ) begin
        s895_val_n7 <= s894_val_n7;
    end
    always @(posedge \clk ) begin
        s895_val_n8 <= s894_val_n8;
    end
    always @(posedge \clk ) begin
        \s896_val  <= \s895_val ;
    end
    always @(posedge \clk ) begin
        s896_val_n1 <= s895_val_n1;
    end
    always @(posedge \clk ) begin
        s896_val_n2 <= s895_val_n2;
    end
    always @(posedge \clk ) begin
        s896_val_n3 <= s895_val_n3;
    end
    always @(posedge \clk ) begin
        s896_val_n4 <= s895_val_n4;
    end
    always @(posedge \clk ) begin
        s896_val_n5 <= s895_val_n5;
    end
    always @(posedge \clk ) begin
        s896_val_n6 <= s895_val_n6;
    end
    always @(posedge \clk ) begin
        s896_val_n7 <= s895_val_n7;
    end
    always @(posedge \clk ) begin
        s896_val_n8 <= s895_val_n8;
    end
    always @(posedge \clk ) begin
        \s897_val  <= \s896_val ;
    end
    always @(posedge \clk ) begin
        s897_val_n1 <= s896_val_n1;
    end
    always @(posedge \clk ) begin
        s897_val_n2 <= s896_val_n2;
    end
    always @(posedge \clk ) begin
        s897_val_n3 <= s896_val_n3;
    end
    always @(posedge \clk ) begin
        s897_val_n4 <= s896_val_n4;
    end
    always @(posedge \clk ) begin
        s897_val_n5 <= s896_val_n5;
    end
    always @(posedge \clk ) begin
        s897_val_n6 <= s896_val_n6;
    end
    always @(posedge \clk ) begin
        s897_val_n7 <= s896_val_n7;
    end
    always @(posedge \clk ) begin
        s897_val_n8 <= s896_val_n8;
    end
    always @(posedge \clk ) begin
        \s898_val  <= \s897_val ;
    end
    always @(posedge \clk ) begin
        s898_val_n1 <= s897_val_n1;
    end
    always @(posedge \clk ) begin
        s898_val_n2 <= s897_val_n2;
    end
    always @(posedge \clk ) begin
        s898_val_n3 <= s897_val_n3;
    end
    always @(posedge \clk ) begin
        s898_val_n4 <= s897_val_n4;
    end
    always @(posedge \clk ) begin
        s898_val_n5 <= s897_val_n5;
    end
    always @(posedge \clk ) begin
        s898_val_n6 <= s897_val_n6;
    end
    always @(posedge \clk ) begin
        s898_val_n7 <= s897_val_n7;
    end
    always @(posedge \clk ) begin
        s898_val_n8 <= s897_val_n8;
    end
    always @(posedge \clk ) begin
        \s899_val  <= \s898_val ;
    end
    always @(posedge \clk ) begin
        s899_val_n1 <= s898_val_n1;
    end
    always @(posedge \clk ) begin
        s899_val_n2 <= s898_val_n2;
    end
    always @(posedge \clk ) begin
        s899_val_n3 <= s898_val_n3;
    end
    always @(posedge \clk ) begin
        s899_val_n4 <= s898_val_n4;
    end
    always @(posedge \clk ) begin
        s899_val_n5 <= s898_val_n5;
    end
    always @(posedge \clk ) begin
        s899_val_n6 <= s898_val_n6;
    end
    always @(posedge \clk ) begin
        s899_val_n7 <= s898_val_n7;
    end
    always @(posedge \clk ) begin
        s899_val_n8 <= s898_val_n8;
    end
    always @(posedge \clk ) begin
        \s900_val  <= \s899_val ;
    end
    always @(posedge \clk ) begin
        s900_val_n1 <= s899_val_n1;
    end
    always @(posedge \clk ) begin
        s900_val_n2 <= s899_val_n2;
    end
    always @(posedge \clk ) begin
        s900_val_n3 <= s899_val_n3;
    end
    always @(posedge \clk ) begin
        s900_val_n4 <= s899_val_n4;
    end
    always @(posedge \clk ) begin
        s900_val_n5 <= s899_val_n5;
    end
    always @(posedge \clk ) begin
        s900_val_n6 <= s899_val_n6;
    end
    always @(posedge \clk ) begin
        s900_val_n7 <= s899_val_n7;
    end
    always @(posedge \clk ) begin
        s900_val_n8 <= s899_val_n8;
    end
    (* src = "src/sreg.spade:127,19" *)
    \tt07_delay_line_tmng::sreg::shift_reg100  shift_reg100_0(.clk_i(\clk ), .val_i(\val ), .output__(val_n1));
    (* src = "src/sreg.spade:129,19" *)
    \tt07_delay_line_tmng::sreg::shift_reg100  shift_reg100_1(.clk_i(\clk ), .val_i(val_n1), .output__(val_n2));
    (* src = "src/sreg.spade:131,19" *)
    \tt07_delay_line_tmng::sreg::shift_reg100  shift_reg100_2(.clk_i(\clk ), .val_i(val_n2), .output__(val_n3));
    (* src = "src/sreg.spade:133,19" *)
    \tt07_delay_line_tmng::sreg::shift_reg100  shift_reg100_3(.clk_i(\clk ), .val_i(val_n3), .output__(val_n4));
    (* src = "src/sreg.spade:135,19" *)
    \tt07_delay_line_tmng::sreg::shift_reg100  shift_reg100_4(.clk_i(\clk ), .val_i(val_n4), .output__(val_n5));
    (* src = "src/sreg.spade:137,19" *)
    \tt07_delay_line_tmng::sreg::shift_reg100  shift_reg100_5(.clk_i(\clk ), .val_i(val_n5), .output__(val_n6));
    (* src = "src/sreg.spade:139,19" *)
    \tt07_delay_line_tmng::sreg::shift_reg100  shift_reg100_6(.clk_i(\clk ), .val_i(val_n6), .output__(val_n7));
    (* src = "src/sreg.spade:141,19" *)
    \tt07_delay_line_tmng::sreg::shift_reg100  shift_reg100_7(.clk_i(\clk ), .val_i(val_n7), .output__(val_n8));
    (* src = "src/sreg.spade:143,19" *)
    \tt07_delay_line_tmng::sreg::shift_reg100  shift_reg100_8(.clk_i(\clk ), .val_i(val_n8), .output__(val_n9));
    assign output__ = val_n9;
endmodule

module \tt07_delay_line_tmng::main::tmng  (
        input clk_i,
        input[5:0] ctrl_i,
        output[7:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "tt07_delay_line_tmng::main::tmng" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \tt07_delay_line_tmng::main::tmng );
        end
    end
    `endif
    logic \clk ;
    assign \clk  = clk_i;
    logic[5:0] \ctrl ;
    assign \ctrl  = ctrl_i;
    (* src = "src/main.spade:16,23" *)
    logic _e_874;
    (* src = "src/main.spade:16,20" *)
    logic _e_873;
    (* src = "src/main.spade:16,14" *)
    reg \opa ;
    (* src = "src/main.spade:17,23" *)
    logic _e_883;
    (* src = "src/main.spade:17,20" *)
    logic _e_882;
    (* src = "src/main.spade:17,14" *)
    reg \opb ;
    (* src = "src/main.spade:18,18" *)
    logic _e_890;
    (* src = "src/main.spade:18,16" *)
    logic \nand ;
    (* src = "src/main.spade:20,22" *)
    logic _e_895;
    (* src = "src/main.spade:22,15" *)
    logic _e_900;
    (* src = "src/main.spade:23,9" *)
    logic _e_903;
    (* src = "src/main.spade:22,12" *)
    logic _e_899;
    (* src = "src/main.spade:20,19" *)
    logic \sreg_in ;
    (* src = "src/main.spade:28,20" *)
    logic \sreg_out ;
    (* src = "src/main.spade:30,33" *)
    logic _e_915;
    logic[7:0] _e_921;
    (* src = "src/main.spade:30,53" *)
    logic[7:0] _e_919;
    logic[7:0] _e_925;
    logic[7:0] _e_927;
    (* src = "src/main.spade:30,75" *)
    logic[7:0] _e_922;
    (* src = "src/main.spade:30,53" *)
    logic[7:0] _e_918;
    (* src = "src/main.spade:30,30" *)
    logic[7:0] _e_914;
    (* src = "src/main.spade:30,14" *)
    reg[7:0] \output_values ;
    assign _e_874 = \ctrl [2];
    assign _e_873 = _e_874 ? \sreg_out  : \opa ;
    always @(posedge \clk ) begin
        \opa  <= _e_873;
    end
    assign _e_883 = \ctrl [1];
    assign _e_882 = _e_883 ? \sreg_out  : \opb ;
    always @(posedge \clk ) begin
        \opb  <= _e_882;
    end
    assign _e_890 = \opa  && \opb ;
    assign \nand  = !_e_890;
    assign _e_895 = \ctrl [5];
    assign _e_900 = \ctrl [4];
    assign _e_903 = \ctrl [3];
    assign _e_899 = _e_900 ? _e_903 : \sreg_out ;
    assign \sreg_in  = _e_895 ? \nand  : _e_899;
    (* src = "src/main.spade:28,20" *)
    \tt07_delay_line_tmng::sreg::shift_reg  shift_reg_0(.clk_i(\clk ), .val_i(\sreg_in ), .output__(\sreg_out ));
    assign _e_915 = \ctrl [0];
    assign _e_921 = 1;
    assign _e_919 = \output_values  << _e_921;
    assign _e_925 = 1;
    assign _e_927 = 0;
    assign _e_922 = \sreg_out  ? _e_925 : _e_927;
    assign _e_918 = _e_919 | _e_922;
    assign _e_914 = _e_915 ? _e_918 : \output_values ;
    always @(posedge \clk ) begin
        \output_values  <= _e_914;
    end
    assign output__ = \output_values ;
endmodule

module tt_um_delay_line_tmng (
        input[7:0] ui_in,
        output[7:0] uo_out,
        input[7:0] uio_in,
        output[7:0] uio_out,
        output[7:0] uio_oe,
        input ena,
        input clk,
        input rst_n
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "tt_um_delay_line_tmng" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, tt_um_delay_line_tmng);
        end
    end
    `endif
    logic[7:0] \uo_out_mut ;
    assign uo_out = \uo_out_mut ;
    logic[7:0] \uio_out_mut ;
    assign uio_out = \uio_out_mut ;
    logic[7:0] \uio_oe_mut ;
    assign uio_oe = \uio_oe_mut ;
    (* src = "src/main.spade:53,14" *)
    reg[7:0] \ui_in_sync ;
    logic[2:0] _e_938;
    (* src = "src/main.spade:56,21" *)
    logic _e_936;
    logic[2:0] _e_941;
    (* src = "src/main.spade:57,22" *)
    logic _e_939;
    logic[2:0] _e_944;
    (* src = "src/main.spade:58,17" *)
    logic _e_942;
    logic[2:0] _e_947;
    (* src = "src/main.spade:59,19" *)
    logic _e_945;
    logic[2:0] _e_950;
    (* src = "src/main.spade:60,19" *)
    logic _e_948;
    logic[2:0] _e_953;
    (* src = "src/main.spade:61,23" *)
    logic _e_951;
    (* src = "src/main.spade:55,16" *)
    logic[5:0] \ctrl ;
    (* src = "src/main.spade:66,18" *)
    logic[7:0] _e_956;
    logic[7:0] _e_960;
    logic[7:0] _e_962;
    always @(posedge \clk ) begin
        \ui_in_sync  <= \ui_in ;
    end
    assign _e_938 = 0;
    assign _e_936 = \ui_in_sync [_e_938];
    assign _e_941 = 1;
    assign _e_939 = \ui_in_sync [_e_941];
    assign _e_944 = 2;
    assign _e_942 = \ui_in_sync [_e_944];
    assign _e_947 = 3;
    assign _e_945 = \ui_in_sync [_e_947];
    assign _e_950 = 4;
    assign _e_948 = \ui_in_sync [_e_950];
    assign _e_953 = 5;
    assign _e_951 = \ui_in_sync [_e_953];
    assign \ctrl  = {_e_936, _e_939, _e_942, _e_945, _e_948, _e_951};
    (* src = "src/main.spade:66,18" *)
    \tt07_delay_line_tmng::main::tmng  tmng_0(.clk_i(\clk ), .ctrl_i(\ctrl ), .output__(_e_956));
    assign \uo_out_mut  = _e_956;
    assign _e_960 = 0;
    assign \uio_out_mut  = _e_960;
    assign _e_962 = 0;
    assign \uio_oe_mut  = _e_962;
endmodule

module \std::cdc::unsafe::sync2[431]  (
        input clk_i,
        input in_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::cdc::unsafe::sync2[431]" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::cdc::unsafe::sync2[431] );
        end
    end
    `endif
    logic \clk ;
    assign \clk  = clk_i;
    logic \in ;
    assign \in  = in_i;
    (* src = "<compiler dir>/stdlib/cdc.spade:20,18" *)
    reg \sync1 ;
    (* src = "<compiler dir>/stdlib/cdc.spade:21,18" *)
    reg \sync2 ;
    always @(posedge \clk ) begin
        \sync1  <= \in ;
    end
    always @(posedge \clk ) begin
        \sync2  <= \sync1 ;
    end
    assign output__ = \sync2 ;
endmodule